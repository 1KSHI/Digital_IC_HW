
module DivRom (
    input wire [9:0] in,
    output wire [11:0] div
);
assign div = div_out;
reg [11:0] div_out;
always @(*) begin
case(in)
0    : div_out = 12'd4095;//2^22
1    : div_out = 12'd4092;
2    : div_out = 12'd4088;
3    : div_out = 12'd4084;
4    : div_out = 12'd4080;
5    : div_out = 12'd4076;
6    : div_out = 12'd4072;
7    : div_out = 12'd4068;
8    : div_out = 12'd4064;
9    : div_out = 12'd4060;
10   : div_out = 12'd4056;
11   : div_out = 12'd4052;
12   : div_out = 12'd4049;
13   : div_out = 12'd4045;
14   : div_out = 12'd4041;
15   : div_out = 12'd4037;
16   : div_out = 12'd4033;
17   : div_out = 12'd4029;
18   : div_out = 12'd4025;
19   : div_out = 12'd4021;
20   : div_out = 12'd4018;
21   : div_out = 12'd4014;
22   : div_out = 12'd4010;
23   : div_out = 12'd4006;
24   : div_out = 12'd4002;
25   : div_out = 12'd3998;
26   : div_out = 12'd3995;
27   : div_out = 12'd3991;
28   : div_out = 12'd3987;
29   : div_out = 12'd3983;
30   : div_out = 12'd3979;
31   : div_out = 12'd3976;
32   : div_out = 12'd3972;
33   : div_out = 12'd3968;
34   : div_out = 12'd3964;
35   : div_out = 12'd3961;
36   : div_out = 12'd3957;
37   : div_out = 12'd3953;
38   : div_out = 12'd3949;
39   : div_out = 12'd3946;
40   : div_out = 12'd3942;
41   : div_out = 12'd3938;
42   : div_out = 12'd3935;
43   : div_out = 12'd3931;
44   : div_out = 12'd3927;
45   : div_out = 12'd3924;
46   : div_out = 12'd3920;
47   : div_out = 12'd3916;
48   : div_out = 12'd3913;
49   : div_out = 12'd3909;
50   : div_out = 12'd3905;
51   : div_out = 12'd3902;
52   : div_out = 12'd3898;
53   : div_out = 12'd3894;
54   : div_out = 12'd3891;
55   : div_out = 12'd3887;
56   : div_out = 12'd3884;
57   : div_out = 12'd3880;
58   : div_out = 12'd3876;
59   : div_out = 12'd3873;
60   : div_out = 12'd3869;
61   : div_out = 12'd3866;
62   : div_out = 12'd3862;
63   : div_out = 12'd3859;
64   : div_out = 12'd3855;
65   : div_out = 12'd3852;
66   : div_out = 12'd3848;
67   : div_out = 12'd3844;
68   : div_out = 12'd3841;
69   : div_out = 12'd3837;
70   : div_out = 12'd3834;
71   : div_out = 12'd3830;
72   : div_out = 12'd3827;
73   : div_out = 12'd3823;
74   : div_out = 12'd3820;
75   : div_out = 12'd3816;
76   : div_out = 12'd3813;
77   : div_out = 12'd3810;
78   : div_out = 12'd3806;
79   : div_out = 12'd3803;
80   : div_out = 12'd3799;
81   : div_out = 12'd3796;
82   : div_out = 12'd3792;
83   : div_out = 12'd3789;
84   : div_out = 12'd3785;
85   : div_out = 12'd3782;
86   : div_out = 12'd3779;
87   : div_out = 12'd3775;
88   : div_out = 12'd3772;
89   : div_out = 12'd3768;
90   : div_out = 12'd3765;
91   : div_out = 12'd3762;
92   : div_out = 12'd3758;
93   : div_out = 12'd3755;
94   : div_out = 12'd3752;
95   : div_out = 12'd3748;
96   : div_out = 12'd3745;
97   : div_out = 12'd3742;
98   : div_out = 12'd3738;
99   : div_out = 12'd3735;
100  : div_out = 12'd3732;
101  : div_out = 12'd3728;
102  : div_out = 12'd3725;
103  : div_out = 12'd3722;
104  : div_out = 12'd3718;
105  : div_out = 12'd3715;
106  : div_out = 12'd3712;
107  : div_out = 12'd3708;
108  : div_out = 12'd3705;
109  : div_out = 12'd3702;
110  : div_out = 12'd3699;
111  : div_out = 12'd3695;
112  : div_out = 12'd3692;
113  : div_out = 12'd3689;
114  : div_out = 12'd3686;
115  : div_out = 12'd3682;
116  : div_out = 12'd3679;
117  : div_out = 12'd3676;
118  : div_out = 12'd3673;
119  : div_out = 12'd3670;
120  : div_out = 12'd3666;
121  : div_out = 12'd3663;
122  : div_out = 12'd3660;
123  : div_out = 12'd3657;
124  : div_out = 12'd3654;
125  : div_out = 12'd3650;
126  : div_out = 12'd3647;
127  : div_out = 12'd3644;
128  : div_out = 12'd3641;
129  : div_out = 12'd3638;
130  : div_out = 12'd3635;
131  : div_out = 12'd3631;
132  : div_out = 12'd3628;
133  : div_out = 12'd3625;
134  : div_out = 12'd3622;
135  : div_out = 12'd3619;
136  : div_out = 12'd3616;
137  : div_out = 12'd3613;
138  : div_out = 12'd3610;
139  : div_out = 12'd3606;
140  : div_out = 12'd3603;
141  : div_out = 12'd3600;
142  : div_out = 12'd3597;
143  : div_out = 12'd3594;
144  : div_out = 12'd3591;
145  : div_out = 12'd3588;
146  : div_out = 12'd3585;
147  : div_out = 12'd3582;
148  : div_out = 12'd3579;
149  : div_out = 12'd3576;
150  : div_out = 12'd3573;
151  : div_out = 12'd3570;
152  : div_out = 12'd3567;
153  : div_out = 12'd3564;
154  : div_out = 12'd3561;
155  : div_out = 12'd3558;
156  : div_out = 12'd3554;
157  : div_out = 12'd3551;
158  : div_out = 12'd3548;
159  : div_out = 12'd3545;
160  : div_out = 12'd3542;
161  : div_out = 12'd3539;
162  : div_out = 12'd3537;
163  : div_out = 12'd3534;
164  : div_out = 12'd3531;
165  : div_out = 12'd3528;
166  : div_out = 12'd3525;
167  : div_out = 12'd3522;
168  : div_out = 12'd3519;
169  : div_out = 12'd3516;
170  : div_out = 12'd3513;
171  : div_out = 12'd3510;
172  : div_out = 12'd3507;
173  : div_out = 12'd3504;
174  : div_out = 12'd3501;
175  : div_out = 12'd3498;
176  : div_out = 12'd3495;
177  : div_out = 12'd3492;
178  : div_out = 12'd3489;
179  : div_out = 12'd3487;
180  : div_out = 12'd3484;
181  : div_out = 12'd3481;
182  : div_out = 12'd3478;
183  : div_out = 12'd3475;
184  : div_out = 12'd3472;
185  : div_out = 12'd3469;
186  : div_out = 12'd3466;
187  : div_out = 12'd3464;
188  : div_out = 12'd3461;
189  : div_out = 12'd3458;
190  : div_out = 12'd3455;
191  : div_out = 12'd3452;
192  : div_out = 12'd3449;
193  : div_out = 12'd3446;
194  : div_out = 12'd3444;
195  : div_out = 12'd3441;
196  : div_out = 12'd3438;
197  : div_out = 12'd3435;
198  : div_out = 12'd3432;
199  : div_out = 12'd3430;
200  : div_out = 12'd3427;
201  : div_out = 12'd3424;
202  : div_out = 12'd3421;
203  : div_out = 12'd3418;
204  : div_out = 12'd3416;
205  : div_out = 12'd3413;
206  : div_out = 12'd3410;
207  : div_out = 12'd3407;
208  : div_out = 12'd3404;
209  : div_out = 12'd3402;
210  : div_out = 12'd3399;
211  : div_out = 12'd3396;
212  : div_out = 12'd3393;
213  : div_out = 12'd3391;
214  : div_out = 12'd3388;
215  : div_out = 12'd3385;
216  : div_out = 12'd3383;
217  : div_out = 12'd3380;
218  : div_out = 12'd3377;
219  : div_out = 12'd3374;
220  : div_out = 12'd3372;
221  : div_out = 12'd3369;
222  : div_out = 12'd3366;
223  : div_out = 12'd3364;
224  : div_out = 12'd3361;
225  : div_out = 12'd3358;
226  : div_out = 12'd3355;
227  : div_out = 12'd3353;
228  : div_out = 12'd3350;
229  : div_out = 12'd3347;
230  : div_out = 12'd3345;
231  : div_out = 12'd3342;
232  : div_out = 12'd3339;
233  : div_out = 12'd3337;
234  : div_out = 12'd3334;
235  : div_out = 12'd3331;
236  : div_out = 12'd3329;
237  : div_out = 12'd3326;
238  : div_out = 12'd3324;
239  : div_out = 12'd3321;
240  : div_out = 12'd3318;
241  : div_out = 12'd3316;
242  : div_out = 12'd3313;
243  : div_out = 12'd3310;
244  : div_out = 12'd3308;
245  : div_out = 12'd3305;
246  : div_out = 12'd3303;
247  : div_out = 12'd3300;
248  : div_out = 12'd3297;
249  : div_out = 12'd3295;
250  : div_out = 12'd3292;
251  : div_out = 12'd3290;
252  : div_out = 12'd3287;
253  : div_out = 12'd3284;
254  : div_out = 12'd3282;
255  : div_out = 12'd3279;
256  : div_out = 12'd3277;
257  : div_out = 12'd3274;
258  : div_out = 12'd3272;
259  : div_out = 12'd3269;
260  : div_out = 12'd3267;
261  : div_out = 12'd3264;
262  : div_out = 12'd3262;
263  : div_out = 12'd3259;
264  : div_out = 12'd3256;
265  : div_out = 12'd3254;
266  : div_out = 12'd3251;
267  : div_out = 12'd3249;
268  : div_out = 12'd3246;
269  : div_out = 12'd3244;
270  : div_out = 12'd3241;
271  : div_out = 12'd3239;
272  : div_out = 12'd3236;
273  : div_out = 12'd3234;
274  : div_out = 12'd3231;
275  : div_out = 12'd3229;
276  : div_out = 12'd3226;
277  : div_out = 12'd3224;
278  : div_out = 12'd3221;
279  : div_out = 12'd3219;
280  : div_out = 12'd3216;
281  : div_out = 12'd3214;
282  : div_out = 12'd3212;
283  : div_out = 12'd3209;
284  : div_out = 12'd3207;
285  : div_out = 12'd3204;
286  : div_out = 12'd3202;
287  : div_out = 12'd3199;
288  : div_out = 12'd3197;
289  : div_out = 12'd3194;
290  : div_out = 12'd3192;
291  : div_out = 12'd3190;
292  : div_out = 12'd3187;
293  : div_out = 12'd3185;
294  : div_out = 12'd3182;
295  : div_out = 12'd3180;
296  : div_out = 12'd3178;
297  : div_out = 12'd3175;
298  : div_out = 12'd3173;
299  : div_out = 12'd3170;
300  : div_out = 12'd3168;
301  : div_out = 12'd3166;
302  : div_out = 12'd3163;
303  : div_out = 12'd3161;
304  : div_out = 12'd3158;
305  : div_out = 12'd3156;
306  : div_out = 12'd3154;
307  : div_out = 12'd3151;
308  : div_out = 12'd3149;
309  : div_out = 12'd3147;
310  : div_out = 12'd3144;
311  : div_out = 12'd3142;
312  : div_out = 12'd3139;
313  : div_out = 12'd3137;
314  : div_out = 12'd3135;
315  : div_out = 12'd3132;
316  : div_out = 12'd3130;
317  : div_out = 12'd3128;
318  : div_out = 12'd3125;
319  : div_out = 12'd3123;
320  : div_out = 12'd3121;
321  : div_out = 12'd3118;
322  : div_out = 12'd3116;
323  : div_out = 12'd3114;
324  : div_out = 12'd3112;
325  : div_out = 12'd3109;
326  : div_out = 12'd3107;
327  : div_out = 12'd3105;
328  : div_out = 12'd3102;
329  : div_out = 12'd3100;
330  : div_out = 12'd3098;
331  : div_out = 12'd3095;
332  : div_out = 12'd3093;
333  : div_out = 12'd3091;
334  : div_out = 12'd3089;
335  : div_out = 12'd3086;
336  : div_out = 12'd3084;
337  : div_out = 12'd3082;
338  : div_out = 12'd3080;
339  : div_out = 12'd3077;
340  : div_out = 12'd3075;
341  : div_out = 12'd3073;
342  : div_out = 12'd3071;
343  : div_out = 12'd3068;
344  : div_out = 12'd3066;
345  : div_out = 12'd3064;
346  : div_out = 12'd3062;
347  : div_out = 12'd3059;
348  : div_out = 12'd3057;
349  : div_out = 12'd3055;
350  : div_out = 12'd3053;
351  : div_out = 12'd3050;
352  : div_out = 12'd3048;
353  : div_out = 12'd3046;
354  : div_out = 12'd3044;
355  : div_out = 12'd3042;
356  : div_out = 12'd3039;
357  : div_out = 12'd3037;
358  : div_out = 12'd3035;
359  : div_out = 12'd3033;
360  : div_out = 12'd3031;
361  : div_out = 12'd3028;
362  : div_out = 12'd3026;
363  : div_out = 12'd3024;
364  : div_out = 12'd3022;
365  : div_out = 12'd3020;
366  : div_out = 12'd3017;
367  : div_out = 12'd3015;
368  : div_out = 12'd3013;
369  : div_out = 12'd3011;
370  : div_out = 12'd3009;
371  : div_out = 12'd3007;
372  : div_out = 12'd3005;
373  : div_out = 12'd3002;
374  : div_out = 12'd3000;
375  : div_out = 12'd2998;
376  : div_out = 12'd2996;
377  : div_out = 12'd2994;
378  : div_out = 12'd2992;
379  : div_out = 12'd2990;
380  : div_out = 12'd2987;
381  : div_out = 12'd2985;
382  : div_out = 12'd2983;
383  : div_out = 12'd2981;
384  : div_out = 12'd2979;
385  : div_out = 12'd2977;
386  : div_out = 12'd2975;
387  : div_out = 12'd2973;
388  : div_out = 12'd2970;
389  : div_out = 12'd2968;
390  : div_out = 12'd2966;
391  : div_out = 12'd2964;
392  : div_out = 12'd2962;
393  : div_out = 12'd2960;
394  : div_out = 12'd2958;
395  : div_out = 12'd2956;
396  : div_out = 12'd2954;
397  : div_out = 12'd2952;
398  : div_out = 12'd2950;
399  : div_out = 12'd2948;
400  : div_out = 12'd2945;
401  : div_out = 12'd2943;
402  : div_out = 12'd2941;
403  : div_out = 12'd2939;
404  : div_out = 12'd2937;
405  : div_out = 12'd2935;
406  : div_out = 12'd2933;
407  : div_out = 12'd2931;
408  : div_out = 12'd2929;
409  : div_out = 12'd2927;
410  : div_out = 12'd2925;
411  : div_out = 12'd2923;
412  : div_out = 12'd2921;
413  : div_out = 12'd2919;
414  : div_out = 12'd2917;
415  : div_out = 12'd2915;
416  : div_out = 12'd2913;
417  : div_out = 12'd2911;
418  : div_out = 12'd2909;
419  : div_out = 12'd2907;
420  : div_out = 12'd2905;
421  : div_out = 12'd2903;
422  : div_out = 12'd2901;
423  : div_out = 12'd2899;
424  : div_out = 12'd2897;
425  : div_out = 12'd2895;
426  : div_out = 12'd2893;
427  : div_out = 12'd2891;
428  : div_out = 12'd2889;
429  : div_out = 12'd2887;
430  : div_out = 12'd2885;
431  : div_out = 12'd2883;
432  : div_out = 12'd2881;
433  : div_out = 12'd2879;
434  : div_out = 12'd2877;
435  : div_out = 12'd2875;
436  : div_out = 12'd2873;
437  : div_out = 12'd2871;
438  : div_out = 12'd2869;
439  : div_out = 12'd2867;
440  : div_out = 12'd2865;
441  : div_out = 12'd2863;
442  : div_out = 12'd2861;
443  : div_out = 12'd2859;
444  : div_out = 12'd2857;
445  : div_out = 12'd2855;
446  : div_out = 12'd2853;
447  : div_out = 12'd2851;
448  : div_out = 12'd2849;
449  : div_out = 12'd2847;
450  : div_out = 12'd2846;
451  : div_out = 12'd2844;
452  : div_out = 12'd2842;
453  : div_out = 12'd2840;
454  : div_out = 12'd2838;
455  : div_out = 12'd2836;
456  : div_out = 12'd2834;
457  : div_out = 12'd2832;
458  : div_out = 12'd2830;
459  : div_out = 12'd2828;
460  : div_out = 12'd2826;
461  : div_out = 12'd2824;
462  : div_out = 12'd2823;
463  : div_out = 12'd2821;
464  : div_out = 12'd2819;
465  : div_out = 12'd2817;
466  : div_out = 12'd2815;
467  : div_out = 12'd2813;
468  : div_out = 12'd2811;
469  : div_out = 12'd2809;
470  : div_out = 12'd2807;
471  : div_out = 12'd2806;
472  : div_out = 12'd2804;
473  : div_out = 12'd2802;
474  : div_out = 12'd2800;
475  : div_out = 12'd2798;
476  : div_out = 12'd2796;
477  : div_out = 12'd2794;
478  : div_out = 12'd2792;
479  : div_out = 12'd2791;
480  : div_out = 12'd2789;
481  : div_out = 12'd2787;
482  : div_out = 12'd2785;
483  : div_out = 12'd2783;
484  : div_out = 12'd2781;
485  : div_out = 12'd2780;
486  : div_out = 12'd2778;
487  : div_out = 12'd2776;
488  : div_out = 12'd2774;
489  : div_out = 12'd2772;
490  : div_out = 12'd2770;
491  : div_out = 12'd2769;
492  : div_out = 12'd2767;
493  : div_out = 12'd2765;
494  : div_out = 12'd2763;
495  : div_out = 12'd2761;
496  : div_out = 12'd2759;
497  : div_out = 12'd2758;
498  : div_out = 12'd2756;
499  : div_out = 12'd2754;
500  : div_out = 12'd2752;
501  : div_out = 12'd2750;
502  : div_out = 12'd2749;
503  : div_out = 12'd2747;
504  : div_out = 12'd2745;
505  : div_out = 12'd2743;
506  : div_out = 12'd2741;
507  : div_out = 12'd2740;
508  : div_out = 12'd2738;
509  : div_out = 12'd2736;
510  : div_out = 12'd2734;
511  : div_out = 12'd2732;
512  : div_out = 12'd2731;
513  : div_out = 12'd2729;
514  : div_out = 12'd2727;
515  : div_out = 12'd2725;
516  : div_out = 12'd2724;
517  : div_out = 12'd2722;
518  : div_out = 12'd2720;
519  : div_out = 12'd2718;
520  : div_out = 12'd2717;
521  : div_out = 12'd2715;
522  : div_out = 12'd2713;
523  : div_out = 12'd2711;
524  : div_out = 12'd2709;
525  : div_out = 12'd2708;
526  : div_out = 12'd2706;
527  : div_out = 12'd2704;
528  : div_out = 12'd2703;
529  : div_out = 12'd2701;
530  : div_out = 12'd2699;
531  : div_out = 12'd2697;
532  : div_out = 12'd2696;
533  : div_out = 12'd2694;
534  : div_out = 12'd2692;
535  : div_out = 12'd2690;
536  : div_out = 12'd2689;
537  : div_out = 12'd2687;
538  : div_out = 12'd2685;
539  : div_out = 12'd2683;
540  : div_out = 12'd2682;
541  : div_out = 12'd2680;
542  : div_out = 12'd2678;
543  : div_out = 12'd2677;
544  : div_out = 12'd2675;
545  : div_out = 12'd2673;
546  : div_out = 12'd2672;
547  : div_out = 12'd2670;
548  : div_out = 12'd2668;
549  : div_out = 12'd2666;
550  : div_out = 12'd2665;
551  : div_out = 12'd2663;
552  : div_out = 12'd2661;
553  : div_out = 12'd2660;
554  : div_out = 12'd2658;
555  : div_out = 12'd2656;
556  : div_out = 12'd2655;
557  : div_out = 12'd2653;
558  : div_out = 12'd2651;
559  : div_out = 12'd2650;
560  : div_out = 12'd2648;
561  : div_out = 12'd2646;
562  : div_out = 12'd2645;
563  : div_out = 12'd2643;
564  : div_out = 12'd2641;
565  : div_out = 12'd2640;
566  : div_out = 12'd2638;
567  : div_out = 12'd2636;
568  : div_out = 12'd2635;
569  : div_out = 12'd2633;
570  : div_out = 12'd2631;
571  : div_out = 12'd2630;
572  : div_out = 12'd2628;
573  : div_out = 12'd2626;
574  : div_out = 12'd2625;
575  : div_out = 12'd2623;
576  : div_out = 12'd2621;
577  : div_out = 12'd2620;
578  : div_out = 12'd2618;
579  : div_out = 12'd2617;
580  : div_out = 12'd2615;
581  : div_out = 12'd2613;
582  : div_out = 12'd2612;
583  : div_out = 12'd2610;
584  : div_out = 12'd2608;
585  : div_out = 12'd2607;
586  : div_out = 12'd2605;
587  : div_out = 12'd2604;
588  : div_out = 12'd2602;
589  : div_out = 12'd2600;
590  : div_out = 12'd2599;
591  : div_out = 12'd2597;
592  : div_out = 12'd2595;
593  : div_out = 12'd2594;
594  : div_out = 12'd2592;
595  : div_out = 12'd2591;
596  : div_out = 12'd2589;
597  : div_out = 12'd2587;
598  : div_out = 12'd2586;
599  : div_out = 12'd2584;
600  : div_out = 12'd2583;
601  : div_out = 12'd2581;
602  : div_out = 12'd2580;
603  : div_out = 12'd2578;
604  : div_out = 12'd2576;
605  : div_out = 12'd2575;
606  : div_out = 12'd2573;
607  : div_out = 12'd2572;
608  : div_out = 12'd2570;
609  : div_out = 12'd2568;
610  : div_out = 12'd2567;
611  : div_out = 12'd2565;
612  : div_out = 12'd2564;
613  : div_out = 12'd2562;
614  : div_out = 12'd2561;
615  : div_out = 12'd2559;
616  : div_out = 12'd2558;
617  : div_out = 12'd2556;
618  : div_out = 12'd2554;
619  : div_out = 12'd2553;
620  : div_out = 12'd2551;
621  : div_out = 12'd2550;
622  : div_out = 12'd2548;
623  : div_out = 12'd2547;
624  : div_out = 12'd2545;
625  : div_out = 12'd2544;
626  : div_out = 12'd2542;
627  : div_out = 12'd2540;
628  : div_out = 12'd2539;
629  : div_out = 12'd2537;
630  : div_out = 12'd2536;
631  : div_out = 12'd2534;
632  : div_out = 12'd2533;
633  : div_out = 12'd2531;
634  : div_out = 12'd2530;
635  : div_out = 12'd2528;
636  : div_out = 12'd2527;
637  : div_out = 12'd2525;
638  : div_out = 12'd2524;
639  : div_out = 12'd2522;
640  : div_out = 12'd2521;
641  : div_out = 12'd2519;
642  : div_out = 12'd2518;
643  : div_out = 12'd2516;
644  : div_out = 12'd2515;
645  : div_out = 12'd2513;
646  : div_out = 12'd2512;
647  : div_out = 12'd2510;
648  : div_out = 12'd2509;
649  : div_out = 12'd2507;
650  : div_out = 12'd2506;
651  : div_out = 12'd2504;
652  : div_out = 12'd2503;
653  : div_out = 12'd2501;
654  : div_out = 12'd2500;
655  : div_out = 12'd2498;
656  : div_out = 12'd2497;
657  : div_out = 12'd2495;
658  : div_out = 12'd2494;
659  : div_out = 12'd2492;
660  : div_out = 12'd2491;
661  : div_out = 12'd2489;
662  : div_out = 12'd2488;
663  : div_out = 12'd2486;
664  : div_out = 12'd2485;
665  : div_out = 12'd2483;
666  : div_out = 12'd2482;
667  : div_out = 12'd2480;
668  : div_out = 12'd2479;
669  : div_out = 12'd2477;
670  : div_out = 12'd2476;
671  : div_out = 12'd2475;
672  : div_out = 12'd2473;
673  : div_out = 12'd2472;
674  : div_out = 12'd2470;
675  : div_out = 12'd2469;
676  : div_out = 12'd2467;
677  : div_out = 12'd2466;
678  : div_out = 12'd2464;
679  : div_out = 12'd2463;
680  : div_out = 12'd2461;
681  : div_out = 12'd2460;
682  : div_out = 12'd2459;
683  : div_out = 12'd2457;
684  : div_out = 12'd2456;
685  : div_out = 12'd2454;
686  : div_out = 12'd2453;
687  : div_out = 12'd2451;
688  : div_out = 12'd2450;
689  : div_out = 12'd2449;
690  : div_out = 12'd2447;
691  : div_out = 12'd2446;
692  : div_out = 12'd2444;
693  : div_out = 12'd2443;
694  : div_out = 12'd2441;
695  : div_out = 12'd2440;
696  : div_out = 12'd2439;
697  : div_out = 12'd2437;
698  : div_out = 12'd2436;
699  : div_out = 12'd2434;
700  : div_out = 12'd2433;
701  : div_out = 12'd2431;
702  : div_out = 12'd2430;
703  : div_out = 12'd2429;
704  : div_out = 12'd2427;
705  : div_out = 12'd2426;
706  : div_out = 12'd2424;
707  : div_out = 12'd2423;
708  : div_out = 12'd2422;
709  : div_out = 12'd2420;
710  : div_out = 12'd2419;
711  : div_out = 12'd2417;
712  : div_out = 12'd2416;
713  : div_out = 12'd2415;
714  : div_out = 12'd2413;
715  : div_out = 12'd2412;
716  : div_out = 12'd2411;
717  : div_out = 12'd2409;
718  : div_out = 12'd2408;
719  : div_out = 12'd2406;
720  : div_out = 12'd2405;
721  : div_out = 12'd2404;
722  : div_out = 12'd2402;
723  : div_out = 12'd2401;
724  : div_out = 12'd2399;
725  : div_out = 12'd2398;
726  : div_out = 12'd2397;
727  : div_out = 12'd2395;
728  : div_out = 12'd2394;
729  : div_out = 12'd2393;
730  : div_out = 12'd2391;
731  : div_out = 12'd2390;
732  : div_out = 12'd2389;
733  : div_out = 12'd2387;
734  : div_out = 12'd2386;
735  : div_out = 12'd2384;
736  : div_out = 12'd2383;
737  : div_out = 12'd2382;
738  : div_out = 12'd2380;
739  : div_out = 12'd2379;
740  : div_out = 12'd2378;
741  : div_out = 12'd2376;
742  : div_out = 12'd2375;
743  : div_out = 12'd2374;
744  : div_out = 12'd2372;
745  : div_out = 12'd2371;
746  : div_out = 12'd2370;
747  : div_out = 12'd2368;
748  : div_out = 12'd2367;
749  : div_out = 12'd2366;
750  : div_out = 12'd2364;
751  : div_out = 12'd2363;
752  : div_out = 12'd2362;
753  : div_out = 12'd2360;
754  : div_out = 12'd2359;
755  : div_out = 12'd2358;
756  : div_out = 12'd2356;
757  : div_out = 12'd2355;
758  : div_out = 12'd2354;
759  : div_out = 12'd2352;
760  : div_out = 12'd2351;
761  : div_out = 12'd2350;
762  : div_out = 12'd2348;
763  : div_out = 12'd2347;
764  : div_out = 12'd2346;
765  : div_out = 12'd2344;
766  : div_out = 12'd2343;
767  : div_out = 12'd2342;
768  : div_out = 12'd2341;
769  : div_out = 12'd2339;
770  : div_out = 12'd2338;
771  : div_out = 12'd2337;
772  : div_out = 12'd2335;
773  : div_out = 12'd2334;
774  : div_out = 12'd2333;
775  : div_out = 12'd2331;
776  : div_out = 12'd2330;
777  : div_out = 12'd2329;
778  : div_out = 12'd2328;
779  : div_out = 12'd2326;
780  : div_out = 12'd2325;
781  : div_out = 12'd2324;
782  : div_out = 12'd2322;
783  : div_out = 12'd2321;
784  : div_out = 12'd2320;
785  : div_out = 12'd2319;
786  : div_out = 12'd2317;
787  : div_out = 12'd2316;
788  : div_out = 12'd2315;
789  : div_out = 12'd2313;
790  : div_out = 12'd2312;
791  : div_out = 12'd2311;
792  : div_out = 12'd2310;
793  : div_out = 12'd2308;
794  : div_out = 12'd2307;
795  : div_out = 12'd2306;
796  : div_out = 12'd2305;
797  : div_out = 12'd2303;
798  : div_out = 12'd2302;
799  : div_out = 12'd2301;
800  : div_out = 12'd2300;
801  : div_out = 12'd2298;
802  : div_out = 12'd2297;
803  : div_out = 12'd2296;
804  : div_out = 12'd2294;
805  : div_out = 12'd2293;
806  : div_out = 12'd2292;
807  : div_out = 12'd2291;
808  : div_out = 12'd2289;
809  : div_out = 12'd2288;
810  : div_out = 12'd2287;
811  : div_out = 12'd2286;
812  : div_out = 12'd2284;
813  : div_out = 12'd2283;
814  : div_out = 12'd2282;
815  : div_out = 12'd2281;
816  : div_out = 12'd2280;
817  : div_out = 12'd2278;
818  : div_out = 12'd2277;
819  : div_out = 12'd2276;
820  : div_out = 12'd2275;
821  : div_out = 12'd2273;
822  : div_out = 12'd2272;
823  : div_out = 12'd2271;
824  : div_out = 12'd2270;
825  : div_out = 12'd2268;
826  : div_out = 12'd2267;
827  : div_out = 12'd2266;
828  : div_out = 12'd2265;
829  : div_out = 12'd2264;
830  : div_out = 12'd2262;
831  : div_out = 12'd2261;
832  : div_out = 12'd2260;
833  : div_out = 12'd2259;
834  : div_out = 12'd2257;
835  : div_out = 12'd2256;
836  : div_out = 12'd2255;
837  : div_out = 12'd2254;
838  : div_out = 12'd2253;
839  : div_out = 12'd2251;
840  : div_out = 12'd2250;
841  : div_out = 12'd2249;
842  : div_out = 12'd2248;
843  : div_out = 12'd2247;
844  : div_out = 12'd2245;
845  : div_out = 12'd2244;
846  : div_out = 12'd2243;
847  : div_out = 12'd2242;
848  : div_out = 12'd2241;
849  : div_out = 12'd2239;
850  : div_out = 12'd2238;
851  : div_out = 12'd2237;
852  : div_out = 12'd2236;
853  : div_out = 12'd2235;
854  : div_out = 12'd2233;
855  : div_out = 12'd2232;
856  : div_out = 12'd2231;
857  : div_out = 12'd2230;
858  : div_out = 12'd2229;
859  : div_out = 12'd2227;
860  : div_out = 12'd2226;
861  : div_out = 12'd2225;
862  : div_out = 12'd2224;
863  : div_out = 12'd2223;
864  : div_out = 12'd2222;
865  : div_out = 12'd2220;
866  : div_out = 12'd2219;
867  : div_out = 12'd2218;
868  : div_out = 12'd2217;
869  : div_out = 12'd2216;
870  : div_out = 12'd2215;
871  : div_out = 12'd2213;
872  : div_out = 12'd2212;
873  : div_out = 12'd2211;
874  : div_out = 12'd2210;
875  : div_out = 12'd2209;
876  : div_out = 12'd2208;
877  : div_out = 12'd2206;
878  : div_out = 12'd2205;
879  : div_out = 12'd2204;
880  : div_out = 12'd2203;
881  : div_out = 12'd2202;
882  : div_out = 12'd2201;
883  : div_out = 12'd2199;
884  : div_out = 12'd2198;
885  : div_out = 12'd2197;
886  : div_out = 12'd2196;
887  : div_out = 12'd2195;
888  : div_out = 12'd2194;
889  : div_out = 12'd2193;
890  : div_out = 12'd2191;
891  : div_out = 12'd2190;
892  : div_out = 12'd2189;
893  : div_out = 12'd2188;
894  : div_out = 12'd2187;
895  : div_out = 12'd2186;
896  : div_out = 12'd2185;
897  : div_out = 12'd2183;
898  : div_out = 12'd2182;
899  : div_out = 12'd2181;
900  : div_out = 12'd2180;
901  : div_out = 12'd2179;
902  : div_out = 12'd2178;
903  : div_out = 12'd2177;
904  : div_out = 12'd2175;
905  : div_out = 12'd2174;
906  : div_out = 12'd2173;
907  : div_out = 12'd2172;
908  : div_out = 12'd2171;
909  : div_out = 12'd2170;
910  : div_out = 12'd2169;
911  : div_out = 12'd2168;
912  : div_out = 12'd2166;
913  : div_out = 12'd2165;
914  : div_out = 12'd2164;
915  : div_out = 12'd2163;
916  : div_out = 12'd2162;
917  : div_out = 12'd2161;
918  : div_out = 12'd2160;
919  : div_out = 12'd2159;
920  : div_out = 12'd2158;
921  : div_out = 12'd2156;
922  : div_out = 12'd2155;
923  : div_out = 12'd2154;
924  : div_out = 12'd2153;
925  : div_out = 12'd2152;
926  : div_out = 12'd2151;
927  : div_out = 12'd2150;
928  : div_out = 12'd2149;
929  : div_out = 12'd2148;
930  : div_out = 12'd2147;
931  : div_out = 12'd2145;
932  : div_out = 12'd2144;
933  : div_out = 12'd2143;
934  : div_out = 12'd2142;
935  : div_out = 12'd2141;
936  : div_out = 12'd2140;
937  : div_out = 12'd2139;
938  : div_out = 12'd2138;
939  : div_out = 12'd2137;
940  : div_out = 12'd2136;
941  : div_out = 12'd2135;
942  : div_out = 12'd2133;
943  : div_out = 12'd2132;
944  : div_out = 12'd2131;
945  : div_out = 12'd2130;
946  : div_out = 12'd2129;
947  : div_out = 12'd2128;
948  : div_out = 12'd2127;
949  : div_out = 12'd2126;
950  : div_out = 12'd2125;
951  : div_out = 12'd2124;
952  : div_out = 12'd2123;
953  : div_out = 12'd2122;
954  : div_out = 12'd2120;
955  : div_out = 12'd2119;
956  : div_out = 12'd2118;
957  : div_out = 12'd2117;
958  : div_out = 12'd2116;
959  : div_out = 12'd2115;
960  : div_out = 12'd2114;
961  : div_out = 12'd2113;
962  : div_out = 12'd2112;
963  : div_out = 12'd2111;
964  : div_out = 12'd2110;
965  : div_out = 12'd2109;
966  : div_out = 12'd2108;
967  : div_out = 12'd2107;
968  : div_out = 12'd2106;
969  : div_out = 12'd2105;
970  : div_out = 12'd2103;
971  : div_out = 12'd2102;
972  : div_out = 12'd2101;
973  : div_out = 12'd2100;
974  : div_out = 12'd2099;
975  : div_out = 12'd2098;
976  : div_out = 12'd2097;
977  : div_out = 12'd2096;
978  : div_out = 12'd2095;
979  : div_out = 12'd2094;
980  : div_out = 12'd2093;
981  : div_out = 12'd2092;
982  : div_out = 12'd2091;
983  : div_out = 12'd2090;
984  : div_out = 12'd2089;
985  : div_out = 12'd2088;
986  : div_out = 12'd2087;
987  : div_out = 12'd2086;
988  : div_out = 12'd2085;
989  : div_out = 12'd2084;
990  : div_out = 12'd2083;
991  : div_out = 12'd2082;
992  : div_out = 12'd2081;
993  : div_out = 12'd2079;
994  : div_out = 12'd2078;
995  : div_out = 12'd2077;
996  : div_out = 12'd2076;
997  : div_out = 12'd2075;
998  : div_out = 12'd2074;
999  : div_out = 12'd2073;
1000 : div_out = 12'd2072;
1001 : div_out = 12'd2071;
1002 : div_out = 12'd2070;
1003 : div_out = 12'd2069;
1004 : div_out = 12'd2068;
1005 : div_out = 12'd2067;
1006 : div_out = 12'd2066;
1007 : div_out = 12'd2065;
1008 : div_out = 12'd2064;
1009 : div_out = 12'd2063;
1010 : div_out = 12'd2062;
1011 : div_out = 12'd2061;
1012 : div_out = 12'd2060;
1013 : div_out = 12'd2059;
1014 : div_out = 12'd2058;
1015 : div_out = 12'd2057;
1016 : div_out = 12'd2056;
1017 : div_out = 12'd2055;
1018 : div_out = 12'd2054;
1019 : div_out = 12'd2053;
1020 : div_out = 12'd2052;
1021 : div_out = 12'd2051;
1022 : div_out = 12'd2050;
1023 : div_out = 12'd2049;
default : div_out = 12'd0;
endcase
end

assign div = div_out;
endmodule
