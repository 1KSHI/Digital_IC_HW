module Rom(
    //input clk,
    input [11:0] x_in,
    output reg[12:0] result_out
);

always @(*) begin
    case(x_in)
    0    : result_out = 13'd4095;
    1    : result_out = 13'd4095;
    2    : result_out = 13'd4095;
    3    : result_out = 13'd4095;
    4    : result_out = 13'd4095;
    5    : result_out = 13'd4095;
    6    : result_out = 13'd4095;
    7    : result_out = 13'd4095;
    8    : result_out = 13'd4095;
    9    : result_out = 13'd4095;
    10   : result_out = 13'd4095;
    11   : result_out = 13'd4094;
    12   : result_out = 13'd4094;
    13   : result_out = 13'd4094;
    14   : result_out = 13'd4094;
    15   : result_out = 13'd4094;
    16   : result_out = 13'd4094;
    17   : result_out = 13'd4094;
    18   : result_out = 13'd4093;
    19   : result_out = 13'd4093;
    20   : result_out = 13'd4093;
    21   : result_out = 13'd4093;
    22   : result_out = 13'd4093;
    23   : result_out = 13'd4092;
    24   : result_out = 13'd4092;
    25   : result_out = 13'd4092;
    26   : result_out = 13'd4092;
    27   : result_out = 13'd4091;
    28   : result_out = 13'd4091;
    29   : result_out = 13'd4091;
    30   : result_out = 13'd4091;
    31   : result_out = 13'd4090;
    32   : result_out = 13'd4090;
    33   : result_out = 13'd4090;
    34   : result_out = 13'd4089;
    35   : result_out = 13'd4089;
    36   : result_out = 13'd4089;
    37   : result_out = 13'd4088;
    38   : result_out = 13'd4088;
    39   : result_out = 13'd4088;
    40   : result_out = 13'd4087;
    41   : result_out = 13'd4087;
    42   : result_out = 13'd4087;
    43   : result_out = 13'd4086;
    44   : result_out = 13'd4086;
    45   : result_out = 13'd4085;
    46   : result_out = 13'd4085;
    47   : result_out = 13'd4084;
    48   : result_out = 13'd4084;
    49   : result_out = 13'd4083;
    50   : result_out = 13'd4083;
    51   : result_out = 13'd4082;
    52   : result_out = 13'd4082;
    53   : result_out = 13'd4081;
    54   : result_out = 13'd4081;
    55   : result_out = 13'd4080;
    56   : result_out = 13'd4080;
    57   : result_out = 13'd4079;
    58   : result_out = 13'd4079;
    59   : result_out = 13'd4078;
    60   : result_out = 13'd4078;
    61   : result_out = 13'd4077;
    62   : result_out = 13'd4076;
    63   : result_out = 13'd4076;
    64   : result_out = 13'd4075;
    65   : result_out = 13'd4075;
    66   : result_out = 13'd4074;
    67   : result_out = 13'd4073;
    68   : result_out = 13'd4073;
    69   : result_out = 13'd4072;
    70   : result_out = 13'd4071;
    71   : result_out = 13'd4071;
    72   : result_out = 13'd4070;
    73   : result_out = 13'd4069;
    74   : result_out = 13'd4069;
    75   : result_out = 13'd4068;
    76   : result_out = 13'd4067;
    77   : result_out = 13'd4066;
    78   : result_out = 13'd4066;
    79   : result_out = 13'd4065;
    80   : result_out = 13'd4064;
    81   : result_out = 13'd4063;
    82   : result_out = 13'd4063;
    83   : result_out = 13'd4062;
    84   : result_out = 13'd4061;
    85   : result_out = 13'd4060;
    86   : result_out = 13'd4059;
    87   : result_out = 13'd4059;
    88   : result_out = 13'd4058;
    89   : result_out = 13'd4057;
    90   : result_out = 13'd4056;
    91   : result_out = 13'd4055;
    92   : result_out = 13'd4054;
    93   : result_out = 13'd4053;
    94   : result_out = 13'd4052;
    95   : result_out = 13'd4052;
    96   : result_out = 13'd4051;
    97   : result_out = 13'd4050;
    98   : result_out = 13'd4049;
    99   : result_out = 13'd4048;
    100  : result_out = 13'd4047; 
    101  : result_out = 13'd4046; 
    102  : result_out = 13'd4045; 
    103  : result_out = 13'd4044; 
    104  : result_out = 13'd4043; 
    105  : result_out = 13'd4042; 
    106  : result_out = 13'd4041; 
    107  : result_out = 13'd4040; 
    108  : result_out = 13'd4039; 
    109  : result_out = 13'd4038; 
    110  : result_out = 13'd4037; 
    111  : result_out = 13'd4036; 
    112  : result_out = 13'd4035; 
    113  : result_out = 13'd4034; 
    114  : result_out = 13'd4033; 
    115  : result_out = 13'd4031; 
    116  : result_out = 13'd4030; 
    117  : result_out = 13'd4029; 
    118  : result_out = 13'd4028; 
    119  : result_out = 13'd4027; 
    120  : result_out = 13'd4026; 
    121  : result_out = 13'd4025; 
    122  : result_out = 13'd4023; 
    123  : result_out = 13'd4022; 
    124  : result_out = 13'd4021; 
    125  : result_out = 13'd4020; 
    126  : result_out = 13'd4019; 
    127  : result_out = 13'd4018; 
    128  : result_out = 13'd4016; 
    129  : result_out = 13'd4015; 
    130  : result_out = 13'd4014; 
    131  : result_out = 13'd4013; 
    132  : result_out = 13'd4011; 
    133  : result_out = 13'd4010; 
    134  : result_out = 13'd4009; 
    135  : result_out = 13'd4007; 
    136  : result_out = 13'd4006; 
    137  : result_out = 13'd4005; 
    138  : result_out = 13'd4004; 
    139  : result_out = 13'd4002; 
    140  : result_out = 13'd4001; 
    141  : result_out = 13'd4000; 
    142  : result_out = 13'd3998; 
    143  : result_out = 13'd3997;
    144  : result_out = 13'd3995;
    145  : result_out = 13'd3994;
    146  : result_out = 13'd3993;
    147  : result_out = 13'd3991;
    148  : result_out = 13'd3990;
    149  : result_out = 13'd3988;
    150  : result_out = 13'd3987;
    151  : result_out = 13'd3986;
    152  : result_out = 13'd3984;
    153  : result_out = 13'd3983;
    154  : result_out = 13'd3981;
    155  : result_out = 13'd3980;
    156  : result_out = 13'd3978;
    157  : result_out = 13'd3977;
    158  : result_out = 13'd3975;
    159  : result_out = 13'd3974;
    160  : result_out = 13'd3972;
    161  : result_out = 13'd3971;
    162  : result_out = 13'd3969;
    163  : result_out = 13'd3968;
    164  : result_out = 13'd3966;
    165  : result_out = 13'd3964;
    166  : result_out = 13'd3963;
    167  : result_out = 13'd3961;
    168  : result_out = 13'd3960;
    169  : result_out = 13'd3958;
    170  : result_out = 13'd3957;
    171  : result_out = 13'd3955;
    172  : result_out = 13'd3953;
    173  : result_out = 13'd3952;
    174  : result_out = 13'd3950;
    175  : result_out = 13'd3948;
    176  : result_out = 13'd3947;
    177  : result_out = 13'd3945;
    178  : result_out = 13'd3943;
    179  : result_out = 13'd3942;
    180  : result_out = 13'd3940;
    181  : result_out = 13'd3938;
    182  : result_out = 13'd3936;
    183  : result_out = 13'd3935;
    184  : result_out = 13'd3933;
    185  : result_out = 13'd3931;
    186  : result_out = 13'd3929;
    187  : result_out = 13'd3928;
    188  : result_out = 13'd3926;
    189  : result_out = 13'd3924;
    190  : result_out = 13'd3922;
    191  : result_out = 13'd3920;
    192  : result_out = 13'd3919;
    193  : result_out = 13'd3917;
    194  : result_out = 13'd3915;
    195  : result_out = 13'd3913;
    196  : result_out = 13'd3911;
    197  : result_out = 13'd3909;
    198  : result_out = 13'd3908;
    199  : result_out = 13'd3906;
    200  : result_out = 13'd3904;
    201  : result_out = 13'd3902;
    202  : result_out = 13'd3900;
    203  : result_out = 13'd3898;
    204  : result_out = 13'd3896;
    205  : result_out = 13'd3894;
    206  : result_out = 13'd3892;
    207  : result_out = 13'd3890;
    208  : result_out = 13'd3888;
    209  : result_out = 13'd3886;
    210  : result_out = 13'd3884;
    211  : result_out = 13'd3882;
    212  : result_out = 13'd3880;
    213  : result_out = 13'd3878;
    214  : result_out = 13'd3876;
    215  : result_out = 13'd3874;
    216  : result_out = 13'd3872;
    217  : result_out = 13'd3870;
    218  : result_out = 13'd3868;
    219  : result_out = 13'd3866;
    220  : result_out = 13'd3864;
    221  : result_out = 13'd3862;
    222  : result_out = 13'd3860;
    223  : result_out = 13'd3858;
    224  : result_out = 13'd3856;
    225  : result_out = 13'd3853;
    226  : result_out = 13'd3851;
    227  : result_out = 13'd3849;
    228  : result_out = 13'd3847;
    229  : result_out = 13'd3845;
    230  : result_out = 13'd3843;
    231  : result_out = 13'd3841;
    232  : result_out = 13'd3838;
    233  : result_out = 13'd3836;
    234  : result_out = 13'd3834;
    235  : result_out = 13'd3832;
    236  : result_out = 13'd3830;
    237  : result_out = 13'd3827;
    238  : result_out = 13'd3825;
    239  : result_out = 13'd3823;
    240  : result_out = 13'd3821;
    241  : result_out = 13'd3818;
    242  : result_out = 13'd3816;
    243  : result_out = 13'd3814;
    244  : result_out = 13'd3811;
    245  : result_out = 13'd3809;
    246  : result_out = 13'd3807;
    247  : result_out = 13'd3804;
    248  : result_out = 13'd3802;
    249  : result_out = 13'd3800;
    250  : result_out = 13'd3797;
    251  : result_out = 13'd3795;
    252  : result_out = 13'd3793;
    253  : result_out = 13'd3790;
    254  : result_out = 13'd3788;
    255  : result_out = 13'd3786;
    256  : result_out = 13'd3783;
    257  : result_out = 13'd3781;
    258  : result_out = 13'd3778;
    259  : result_out = 13'd3776;
    260  : result_out = 13'd3774;
    261  : result_out = 13'd3771;
    262  : result_out = 13'd3769;
    263  : result_out = 13'd3766;
    264  : result_out = 13'd3764;
    265  : result_out = 13'd3761;
    266  : result_out = 13'd3759;
    267  : result_out = 13'd3756;
    268  : result_out = 13'd3754;
    269  : result_out = 13'd3751;
    270  : result_out = 13'd3749;
    271  : result_out = 13'd3746;
    272  : result_out = 13'd3744;
    273  : result_out = 13'd3741;
    274  : result_out = 13'd3738;
    275  : result_out = 13'd3736;
    276  : result_out = 13'd3733;
    277  : result_out = 13'd3731;
    278  : result_out = 13'd3728;
    279  : result_out = 13'd3726;
    280  : result_out = 13'd3723;
    281  : result_out = 13'd3720;
    282  : result_out = 13'd3718;
    283  : result_out = 13'd3715;
    284  : result_out = 13'd3712;
    285  : result_out = 13'd3710;
    286  : result_out = 13'd3707;
    287  : result_out = 13'd3704;
    288  : result_out = 13'd3702;
    289  : result_out = 13'd3699;
    290  : result_out = 13'd3696;
    291  : result_out = 13'd3694;
    292  : result_out = 13'd3691;
    293  : result_out = 13'd3688;
    294  : result_out = 13'd3685;
    295  : result_out = 13'd3683;
    296  : result_out = 13'd3680;
    297  : result_out = 13'd3677;
    298  : result_out = 13'd3674;
    299  : result_out = 13'd3672;
    300  : result_out = 13'd3669;
    301  : result_out = 13'd3666;
    302  : result_out = 13'd3663;
    303  : result_out = 13'd3660;
    304  : result_out = 13'd3658;
    305  : result_out = 13'd3655;
    306  : result_out = 13'd3652;
    307  : result_out = 13'd3649;
    308  : result_out = 13'd3646;
    309  : result_out = 13'd3643;
    310  : result_out = 13'd3641;
    311  : result_out = 13'd3638;
    312  : result_out = 13'd3635;
    313  : result_out = 13'd3632;
    314  : result_out = 13'd3629;
    315  : result_out = 13'd3626;
    316  : result_out = 13'd3623;
    317  : result_out = 13'd3620;
    318  : result_out = 13'd3617;
    319  : result_out = 13'd3614;
    320  : result_out = 13'd3611;
    321  : result_out = 13'd3608;
    322  : result_out = 13'd3605;
    323  : result_out = 13'd3602;
    324  : result_out = 13'd3599;
    325  : result_out = 13'd3596;
    326  : result_out = 13'd3593;
    327  : result_out = 13'd3590;
    328  : result_out = 13'd3587;
    329  : result_out = 13'd3584;
    330  : result_out = 13'd3581;
    331  : result_out = 13'd3578;
    332  : result_out = 13'd3575;
    333  : result_out = 13'd3572;
    334  : result_out = 13'd3569;
    335  : result_out = 13'd3566;
    336  : result_out = 13'd3563;
    337  : result_out = 13'd3560;
    338  : result_out = 13'd3557;
    339  : result_out = 13'd3554;
    340  : result_out = 13'd3550;
    341  : result_out = 13'd3547;
    342  : result_out = 13'd3544;
    343  : result_out = 13'd3541;
    344  : result_out = 13'd3538;
    345  : result_out = 13'd3535;
    346  : result_out = 13'd3531;
    347  : result_out = 13'd3528;
    348  : result_out = 13'd3525;
    349  : result_out = 13'd3522;
    350  : result_out = 13'd3519;
    351  : result_out = 13'd3515;
    352  : result_out = 13'd3512;
    353  : result_out = 13'd3509;
    354  : result_out = 13'd3506;
    355  : result_out = 13'd3503;
    356  : result_out = 13'd3499;
    357  : result_out = 13'd3496;
    358  : result_out = 13'd3493;
    359  : result_out = 13'd3489;
    360  : result_out = 13'd3486;
    361  : result_out = 13'd3483;
    362  : result_out = 13'd3480;
    363  : result_out = 13'd3476;
    364  : result_out = 13'd3473;
    365  : result_out = 13'd3470;
    366  : result_out = 13'd3466;
    367  : result_out = 13'd3463;
    368  : result_out = 13'd3460;
    369  : result_out = 13'd3456;
    370  : result_out = 13'd3453;
    371  : result_out = 13'd3449;
    372  : result_out = 13'd3446;
    373  : result_out = 13'd3443;
    374  : result_out = 13'd3439;
    375  : result_out = 13'd3436;
    376  : result_out = 13'd3432;
    377  : result_out = 13'd3429;
    378  : result_out = 13'd3425;
    379  : result_out = 13'd3422;
    380  : result_out = 13'd3419;
    381  : result_out = 13'd3415;
    382  : result_out = 13'd3412;
    383  : result_out = 13'd3408;
    384  : result_out = 13'd3405;
    385  : result_out = 13'd3401;
    386  : result_out = 13'd3398;
    387  : result_out = 13'd3394;
    388  : result_out = 13'd3391;
    389  : result_out = 13'd3387;
    390  : result_out = 13'd3384;
    391  : result_out = 13'd3380;
    392  : result_out = 13'd3377;
    393  : result_out = 13'd3373;
    394  : result_out = 13'd3369;
    395  : result_out = 13'd3366;
    396  : result_out = 13'd3362;
    397  : result_out = 13'd3359;
    398  : result_out = 13'd3355;
    399  : result_out = 13'd3351;
    400  : result_out = 13'd3348;
    401  : result_out = 13'd3344;
    402  : result_out = 13'd3341;
    403  : result_out = 13'd3337;
    404  : result_out = 13'd3333;
    405  : result_out = 13'd3330;
    406  : result_out = 13'd3326;
    407  : result_out = 13'd3322;
    408  : result_out = 13'd3319;
    409  : result_out = 13'd3315;
    410  : result_out = 13'd3311;
    411  : result_out = 13'd3308;
    412  : result_out = 13'd3304;
    413  : result_out = 13'd3300;
    414  : result_out = 13'd3296;
    415  : result_out = 13'd3293;
    416  : result_out = 13'd3289;
    417  : result_out = 13'd3285;
    418  : result_out = 13'd3281;
    419  : result_out = 13'd3278;
    420  : result_out = 13'd3274;
    421  : result_out = 13'd3270;
    422  : result_out = 13'd3266;
    423  : result_out = 13'd3263;
    424  : result_out = 13'd3259;
    425  : result_out = 13'd3255;
    426  : result_out = 13'd3251;
    427  : result_out = 13'd3247;
    428  : result_out = 13'd3243;
    429  : result_out = 13'd3240;
    430  : result_out = 13'd3236;
    431  : result_out = 13'd3232;
    432  : result_out = 13'd3228;
    433  : result_out = 13'd3224;
    434  : result_out = 13'd3220;
    435  : result_out = 13'd3216;
    436  : result_out = 13'd3213;
    437  : result_out = 13'd3209;
    438  : result_out = 13'd3205;
    439  : result_out = 13'd3201;
    440  : result_out = 13'd3197;
    441  : result_out = 13'd3193;
    442  : result_out = 13'd3189;
    443  : result_out = 13'd3185;
    444  : result_out = 13'd3181;
    445  : result_out = 13'd3177;
    446  : result_out = 13'd3173;
    447  : result_out = 13'd3169;
    448  : result_out = 13'd3165;
    449  : result_out = 13'd3161;
    450  : result_out = 13'd3157;
    451  : result_out = 13'd3153;
    452  : result_out = 13'd3149;
    453  : result_out = 13'd3145;
    454  : result_out = 13'd3141;
    455  : result_out = 13'd3137;
    456  : result_out = 13'd3133;
    457  : result_out = 13'd3129;
    458  : result_out = 13'd3125;
    459  : result_out = 13'd3121;
    460  : result_out = 13'd3117;
    461  : result_out = 13'd3113;
    462  : result_out = 13'd3109;
    463  : result_out = 13'd3105;
    464  : result_out = 13'd3101;
    465  : result_out = 13'd3096;
    466  : result_out = 13'd3092;
    467  : result_out = 13'd3088;
    468  : result_out = 13'd3084;
    469  : result_out = 13'd3080;
    470  : result_out = 13'd3076;
    471  : result_out = 13'd3072;
    472  : result_out = 13'd3067;
    473  : result_out = 13'd3063;
    474  : result_out = 13'd3059;
    475  : result_out = 13'd3055;
    476  : result_out = 13'd3051;
    477  : result_out = 13'd3047;
    478  : result_out = 13'd3042;
    479  : result_out = 13'd3038;
    480  : result_out = 13'd3034;
    481  : result_out = 13'd3030;
    482  : result_out = 13'd3025;
    483  : result_out = 13'd3021;
    484  : result_out = 13'd3017;
    485  : result_out = 13'd3013;
    486  : result_out = 13'd3008;
    487  : result_out = 13'd3004;
    488  : result_out = 13'd3000;
    489  : result_out = 13'd2996;
    490  : result_out = 13'd2991;
    491  : result_out = 13'd2987;
    492  : result_out = 13'd2983;
    493  : result_out = 13'd2978;
    494  : result_out = 13'd2974;
    495  : result_out = 13'd2970;
    496  : result_out = 13'd2966;
    497  : result_out = 13'd2961;
    498  : result_out = 13'd2957;
    499  : result_out = 13'd2952;
    500  : result_out = 13'd2948;
    501  : result_out = 13'd2944;
    502  : result_out = 13'd2939;
    503  : result_out = 13'd2935;
    504  : result_out = 13'd2931;
    505  : result_out = 13'd2926;
    506  : result_out = 13'd2922;
    507  : result_out = 13'd2917;
    508  : result_out = 13'd2913;
    509  : result_out = 13'd2909;
    510  : result_out = 13'd2904;
    511  : result_out = 13'd2900;
    512  : result_out = 13'd2895;
    513  : result_out = 13'd2891;
    514  : result_out = 13'd2886;
    515  : result_out = 13'd2882;
    516  : result_out = 13'd2877;
    517  : result_out = 13'd2873;
    518  : result_out = 13'd2869;
    519  : result_out = 13'd2864;
    520  : result_out = 13'd2860;
    521  : result_out = 13'd2855;
    522  : result_out = 13'd2851;
    523  : result_out = 13'd2846;
    524  : result_out = 13'd2842;
    525  : result_out = 13'd2837;
    526  : result_out = 13'd2832;
    527  : result_out = 13'd2828;
    528  : result_out = 13'd2823;
    529  : result_out = 13'd2819;
    530  : result_out = 13'd2814;
    531  : result_out = 13'd2810;
    532  : result_out = 13'd2805;
    533  : result_out = 13'd2801;
    534  : result_out = 13'd2796;
    535  : result_out = 13'd2791;
    536  : result_out = 13'd2787;
    537  : result_out = 13'd2782;
    538  : result_out = 13'd2778;
    539  : result_out = 13'd2773;
    540  : result_out = 13'd2768;
    541  : result_out = 13'd2764;
    542  : result_out = 13'd2759;
    543  : result_out = 13'd2754;
    544  : result_out = 13'd2750;
    545  : result_out = 13'd2745;
    546  : result_out = 13'd2740;
    547  : result_out = 13'd2736;
    548  : result_out = 13'd2731;
    549  : result_out = 13'd2726;
    550  : result_out = 13'd2722;
    551  : result_out = 13'd2717;
    552  : result_out = 13'd2712;
    553  : result_out = 13'd2708;
    554  : result_out = 13'd2703;
    555  : result_out = 13'd2698;
    556  : result_out = 13'd2693;
    557  : result_out = 13'd2689;
    558  : result_out = 13'd2684;
    559  : result_out = 13'd2679;
    560  : result_out = 13'd2674;
    561  : result_out = 13'd2670;
    562  : result_out = 13'd2665;
    563  : result_out = 13'd2660;
    564  : result_out = 13'd2655;
    565  : result_out = 13'd2651;
    566  : result_out = 13'd2646;
    567  : result_out = 13'd2641;
    568  : result_out = 13'd2636;
    569  : result_out = 13'd2631;
    570  : result_out = 13'd2627;
    571  : result_out = 13'd2622;
    572  : result_out = 13'd2617;
    573  : result_out = 13'd2612;
    574  : result_out = 13'd2607;
    575  : result_out = 13'd2602;
    576  : result_out = 13'd2597;
    577  : result_out = 13'd2593;
    578  : result_out = 13'd2588;
    579  : result_out = 13'd2583;
    580  : result_out = 13'd2578;
    581  : result_out = 13'd2573;
    582  : result_out = 13'd2568;
    583  : result_out = 13'd2563;
    584  : result_out = 13'd2558;
    585  : result_out = 13'd2554;
    586  : result_out = 13'd2549;
    587  : result_out = 13'd2544;
    588  : result_out = 13'd2539;
    589  : result_out = 13'd2534;
    590  : result_out = 13'd2529;
    591  : result_out = 13'd2524;
    592  : result_out = 13'd2519;
    593  : result_out = 13'd2514;
    594  : result_out = 13'd2509;
    595  : result_out = 13'd2504;
    596  : result_out = 13'd2499;
    597  : result_out = 13'd2494;
    598  : result_out = 13'd2489;
    599  : result_out = 13'd2484;
    600  : result_out = 13'd2479;
    601  : result_out = 13'd2474;
    602  : result_out = 13'd2469;
    603  : result_out = 13'd2464;
    604  : result_out = 13'd2459;
    605  : result_out = 13'd2454;
    606  : result_out = 13'd2449;
    607  : result_out = 13'd2444;
    608  : result_out = 13'd2439;
    609  : result_out = 13'd2434;
    610  : result_out = 13'd2429;
    611  : result_out = 13'd2424;
    612  : result_out = 13'd2419;
    613  : result_out = 13'd2414;
    614  : result_out = 13'd2409;
    615  : result_out = 13'd2404;
    616  : result_out = 13'd2398;
    617  : result_out = 13'd2393;
    618  : result_out = 13'd2388;
    619  : result_out = 13'd2383;
    620  : result_out = 13'd2378;
    621  : result_out = 13'd2373;
    622  : result_out = 13'd2368;
    623  : result_out = 13'd2363;
    624  : result_out = 13'd2358;
    625  : result_out = 13'd2352;
    626  : result_out = 13'd2347;
    627  : result_out = 13'd2342;
    628  : result_out = 13'd2337;
    629  : result_out = 13'd2332;
    630  : result_out = 13'd2327;
    631  : result_out = 13'd2321;
    632  : result_out = 13'd2316;
    633  : result_out = 13'd2311;
    634  : result_out = 13'd2306;
    635  : result_out = 13'd2301;
    636  : result_out = 13'd2295;
    637  : result_out = 13'd2290;
    638  : result_out = 13'd2285;
    639  : result_out = 13'd2280;
    640  : result_out = 13'd2275;
    641  : result_out = 13'd2269;
    642  : result_out = 13'd2264;
    643  : result_out = 13'd2259;
    644  : result_out = 13'd2254;
    645  : result_out = 13'd2248;
    646  : result_out = 13'd2243;
    647  : result_out = 13'd2238;
    648  : result_out = 13'd2233;
    649  : result_out = 13'd2227;
    650  : result_out = 13'd2222;
    651  : result_out = 13'd2217;
    652  : result_out = 13'd2212;
    653  : result_out = 13'd2206;
    654  : result_out = 13'd2201;
    655  : result_out = 13'd2196;
    656  : result_out = 13'd2190;
    657  : result_out = 13'd2185;
    658  : result_out = 13'd2180;
    659  : result_out = 13'd2174;
    660  : result_out = 13'd2169;
    661  : result_out = 13'd2164;
    662  : result_out = 13'd2158;
    663  : result_out = 13'd2153;
    664  : result_out = 13'd2148;
    665  : result_out = 13'd2142;
    666  : result_out = 13'd2137;
    667  : result_out = 13'd2132;
    668  : result_out = 13'd2126;
    669  : result_out = 13'd2121;
    670  : result_out = 13'd2116;
    671  : result_out = 13'd2110;
    672  : result_out = 13'd2105;
    673  : result_out = 13'd2099;
    674  : result_out = 13'd2094;
    675  : result_out = 13'd2089;
    676  : result_out = 13'd2083;
    677  : result_out = 13'd2078;
    678  : result_out = 13'd2072;
    679  : result_out = 13'd2067;
    680  : result_out = 13'd2061;
    681  : result_out = 13'd2056;
    682  : result_out = 13'd2051;
    683  : result_out = 13'd2045;
    684  : result_out = 13'd2040;
    685  : result_out = 13'd2034;
    686  : result_out = 13'd2029;
    687  : result_out = 13'd2023;
    688  : result_out = 13'd2018;
    689  : result_out = 13'd2012;
    690  : result_out = 13'd2007;
    691  : result_out = 13'd2001;
    692  : result_out = 13'd1996;
    693  : result_out = 13'd1991;
    694  : result_out = 13'd1985;
    695  : result_out = 13'd1980;
    696  : result_out = 13'd1974;
    697  : result_out = 13'd1969;
    698  : result_out = 13'd1963;
    699  : result_out = 13'd1957;
    700  : result_out = 13'd1952;
    701  : result_out = 13'd1946;
    702  : result_out = 13'd1941;
    703  : result_out = 13'd1935;
    704  : result_out = 13'd1930;
    705  : result_out = 13'd1924;
    706  : result_out = 13'd1919;
    707  : result_out = 13'd1913;
    708  : result_out = 13'd1908;
    709  : result_out = 13'd1902;
    710  : result_out = 13'd1897;
    711  : result_out = 13'd1891;
    712  : result_out = 13'd1885;
    713  : result_out = 13'd1880;
    714  : result_out = 13'd1874;
    715  : result_out = 13'd1869;
    716  : result_out = 13'd1863;
    717  : result_out = 13'd1857;
    718  : result_out = 13'd1852;
    719  : result_out = 13'd1846;
    720  : result_out = 13'd1841;
    721  : result_out = 13'd1835;
    722  : result_out = 13'd1829;
    723  : result_out = 13'd1824;
    724  : result_out = 13'd1818;
    725  : result_out = 13'd1812;
    726  : result_out = 13'd1807;
    727  : result_out = 13'd1801;
    728  : result_out = 13'd1796;
    729  : result_out = 13'd1790;
    730  : result_out = 13'd1784;
    731  : result_out = 13'd1779;
    732  : result_out = 13'd1773;
    733  : result_out = 13'd1767;
    734  : result_out = 13'd1762;
    735  : result_out = 13'd1756;
    736  : result_out = 13'd1750;
    737  : result_out = 13'd1745;
    738  : result_out = 13'd1739;
    739  : result_out = 13'd1733;
    740  : result_out = 13'd1728;
    741  : result_out = 13'd1722;
    742  : result_out = 13'd1716;
    743  : result_out = 13'd1710;
    744  : result_out = 13'd1705;
    745  : result_out = 13'd1699;
    746  : result_out = 13'd1693;
    747  : result_out = 13'd1688;
    748  : result_out = 13'd1682;
    749  : result_out = 13'd1676;
    750  : result_out = 13'd1670;
    751  : result_out = 13'd1665;
    752  : result_out = 13'd1659;
    753  : result_out = 13'd1653;
    754  : result_out = 13'd1647;
    755  : result_out = 13'd1642;
    756  : result_out = 13'd1636;
    757  : result_out = 13'd1630;
    758  : result_out = 13'd1624;
    759  : result_out = 13'd1619;
    760  : result_out = 13'd1613;
    761  : result_out = 13'd1607;
    762  : result_out = 13'd1601;
    763  : result_out = 13'd1595;
    764  : result_out = 13'd1590;
    765  : result_out = 13'd1584;
    766  : result_out = 13'd1578;
    767  : result_out = 13'd1572;
    768  : result_out = 13'd1566;
    769  : result_out = 13'd1561;
    770  : result_out = 13'd1555;
    771  : result_out = 13'd1549;
    772  : result_out = 13'd1543;
    773  : result_out = 13'd1537;
    774  : result_out = 13'd1532;
    775  : result_out = 13'd1526;
    776  : result_out = 13'd1520;
    777  : result_out = 13'd1514;
    778  : result_out = 13'd1508;
    779  : result_out = 13'd1502;
    780  : result_out = 13'd1497;
    781  : result_out = 13'd1491;
    782  : result_out = 13'd1485;
    783  : result_out = 13'd1479;
    784  : result_out = 13'd1473;
    785  : result_out = 13'd1467;
    786  : result_out = 13'd1461;
    787  : result_out = 13'd1456;
    788  : result_out = 13'd1450;
    789  : result_out = 13'd1444;
    790  : result_out = 13'd1438;
    791  : result_out = 13'd1432;
    792  : result_out = 13'd1426;
    793  : result_out = 13'd1420;
    794  : result_out = 13'd1414;
    795  : result_out = 13'd1408;
    796  : result_out = 13'd1403;
    797  : result_out = 13'd1397;
    798  : result_out = 13'd1391;
    799  : result_out = 13'd1385;
    800  : result_out = 13'd1379;
    801  : result_out = 13'd1373;
    802  : result_out = 13'd1367;
    803  : result_out = 13'd1361;
    804  : result_out = 13'd1355;
    805  : result_out = 13'd1349;
    806  : result_out = 13'd1343;
    807  : result_out = 13'd1337;
    808  : result_out = 13'd1331;
    809  : result_out = 13'd1326;
    810  : result_out = 13'd1320;
    811  : result_out = 13'd1314;
    812  : result_out = 13'd1308;
    813  : result_out = 13'd1302;
    814  : result_out = 13'd1296;
    815  : result_out = 13'd1290;
    816  : result_out = 13'd1284;
    817  : result_out = 13'd1278;
    818  : result_out = 13'd1272;
    819  : result_out = 13'd1266;
    820  : result_out = 13'd1260;
    821  : result_out = 13'd1254;
    822  : result_out = 13'd1248;
    823  : result_out = 13'd1242;
    824  : result_out = 13'd1236;
    825  : result_out = 13'd1230;
    826  : result_out = 13'd1224;
    827  : result_out = 13'd1218;
    828  : result_out = 13'd1212;
    829  : result_out = 13'd1206;
    830  : result_out = 13'd1200;
    831  : result_out = 13'd1194;
    832  : result_out = 13'd1188;
    833  : result_out = 13'd1182;
    834  : result_out = 13'd1176;
    835  : result_out = 13'd1170;
    836  : result_out = 13'd1164;
    837  : result_out = 13'd1158;
    838  : result_out = 13'd1152;
    839  : result_out = 13'd1146;
    840  : result_out = 13'd1140;
    841  : result_out = 13'd1134;
    842  : result_out = 13'd1128;
    843  : result_out = 13'd1122;
    844  : result_out = 13'd1116;
    845  : result_out = 13'd1110;
    846  : result_out = 13'd1104;
    847  : result_out = 13'd1098;
    848  : result_out = 13'd1091;
    849  : result_out = 13'd1085;
    850  : result_out = 13'd1079;
    851  : result_out = 13'd1073;
    852  : result_out = 13'd1067;
    853  : result_out = 13'd1061;
    854  : result_out = 13'd1055;
    855  : result_out = 13'd1049;
    856  : result_out = 13'd1043;
    857  : result_out = 13'd1037;
    858  : result_out = 13'd1031;
    859  : result_out = 13'd1025;
    860  : result_out = 13'd1019;
    861  : result_out = 13'd1013;
    862  : result_out = 13'd1006;
    863  : result_out = 13'd1000;
    864  : result_out = 13'd994;
    865  : result_out = 13'd988;
    866  : result_out = 13'd982;
    867  : result_out = 13'd976;
    868  : result_out = 13'd970;
    869  : result_out = 13'd964;
    870  : result_out = 13'd958;
    871  : result_out = 13'd952;
    872  : result_out = 13'd945;
    873  : result_out = 13'd939;
    874  : result_out = 13'd933;
    875  : result_out = 13'd927;
    876  : result_out = 13'd921;
    877  : result_out = 13'd915;
    878  : result_out = 13'd909;
    879  : result_out = 13'd903;
    880  : result_out = 13'd896;
    881  : result_out = 13'd890;
    882  : result_out = 13'd884;
    883  : result_out = 13'd878;
    884  : result_out = 13'd872;
    885  : result_out = 13'd866;
    886  : result_out = 13'd860;
    887  : result_out = 13'd853;
    888  : result_out = 13'd847;
    889  : result_out = 13'd841;
    890  : result_out = 13'd835;
    891  : result_out = 13'd829;
    892  : result_out = 13'd823;
    893  : result_out = 13'd817;
    894  : result_out = 13'd810;
    895  : result_out = 13'd804;
    896  : result_out = 13'd798;
    897  : result_out = 13'd792;
    898  : result_out = 13'd786;
    899  : result_out = 13'd780;
    900  : result_out = 13'd773;
    901  : result_out = 13'd767;
    902  : result_out = 13'd761;
    903  : result_out = 13'd755;
    904  : result_out = 13'd749;
    905  : result_out = 13'd743;
    906  : result_out = 13'd736;
    907  : result_out = 13'd730;
    908  : result_out = 13'd724;
    909  : result_out = 13'd718;
    910  : result_out = 13'd712;
    911  : result_out = 13'd705;
    912  : result_out = 13'd699;
    913  : result_out = 13'd693;
    914  : result_out = 13'd687;
    915  : result_out = 13'd681;
    916  : result_out = 13'd674;
    917  : result_out = 13'd668;
    918  : result_out = 13'd662;
    919  : result_out = 13'd656;
    920  : result_out = 13'd650;
    921  : result_out = 13'd643;
    922  : result_out = 13'd637;
    923  : result_out = 13'd631;
    924  : result_out = 13'd625;
    925  : result_out = 13'd619;
    926  : result_out = 13'd612;
    927  : result_out = 13'd606;
    928  : result_out = 13'd600;
    929  : result_out = 13'd594;
    930  : result_out = 13'd588;
    931  : result_out = 13'd581;
    932  : result_out = 13'd575;
    933  : result_out = 13'd569;
    934  : result_out = 13'd563;
    935  : result_out = 13'd556;
    936  : result_out = 13'd550;
    937  : result_out = 13'd544;
    938  : result_out = 13'd538;
    939  : result_out = 13'd532;
    940  : result_out = 13'd525;
    941  : result_out = 13'd519;
    942  : result_out = 13'd513;
    943  : result_out = 13'd507;
    944  : result_out = 13'd500;
    945  : result_out = 13'd494;
    946  : result_out = 13'd488;
    947  : result_out = 13'd482;
    948  : result_out = 13'd475;
    949  : result_out = 13'd469;
    950  : result_out = 13'd463;
    951  : result_out = 13'd457;
    952  : result_out = 13'd450;
    953  : result_out = 13'd444;
    954  : result_out = 13'd438;
    955  : result_out = 13'd432;
    956  : result_out = 13'd425;
    957  : result_out = 13'd419;
    958  : result_out = 13'd413;
    959  : result_out = 13'd407;
    960  : result_out = 13'd400;
    961  : result_out = 13'd394;
    962  : result_out = 13'd388;
    963  : result_out = 13'd382;
    964  : result_out = 13'd375;
    965  : result_out = 13'd369;
    966  : result_out = 13'd363;
    967  : result_out = 13'd357;
    968  : result_out = 13'd350;
    969  : result_out = 13'd344;
    970  : result_out = 13'd338;
    971  : result_out = 13'd332;
    972  : result_out = 13'd325;
    973  : result_out = 13'd319;
    974  : result_out = 13'd313;
    975  : result_out = 13'd307;
    976  : result_out = 13'd300;
    977  : result_out = 13'd294;
    978  : result_out = 13'd288;
    979  : result_out = 13'd282;
    980  : result_out = 13'd275;
    981  : result_out = 13'd269;
    982  : result_out = 13'd263;
    983  : result_out = 13'd256;
    984  : result_out = 13'd250;
    985  : result_out = 13'd244;
    986  : result_out = 13'd238;
    987  : result_out = 13'd231;
    988  : result_out = 13'd225;
    989  : result_out = 13'd219;
    990  : result_out = 13'd213;
    991  : result_out = 13'd206;
    992  : result_out = 13'd200;
    993  : result_out = 13'd194;
    994  : result_out = 13'd187;
    995  : result_out = 13'd181;
    996  : result_out = 13'd175;
    997  : result_out = 13'd169;
    998  : result_out = 13'd162;
    999  : result_out = 13'd156;
    1000 : result_out = 13'd150;
    1001 : result_out = 13'd143;
    1002 : result_out = 13'd137;
    1003 : result_out = 13'd131;
    1004 : result_out = 13'd125;
    1005 : result_out = 13'd118;
    1006 : result_out = 13'd112;
    1007 : result_out = 13'd106;
    1008 : result_out = 13'd100;
    1009 : result_out = 13'd93;
    1010 : result_out = 13'd87;
    1011 : result_out = 13'd81;
    1012 : result_out = 13'd74;
    1013 : result_out = 13'd68;
    1014 : result_out = 13'd62;
    1015 : result_out = 13'd56;
    1016 : result_out = 13'd49;
    1017 : result_out = 13'd43;
    1018 : result_out = 13'd37;
    1019 : result_out = 13'd30;
    1020 : result_out = 13'd24;
    1021 : result_out = 13'd18;
    1022 : result_out = 13'd12;
    1023 : result_out = 13'd5;
    1024 : result_out = 13'd0;
    1025 : result_out = {1'b1,12'd5   };
    1026 : result_out = {1'b1,12'd12  };
    1027 : result_out = {1'b1,12'd18  };
    1028 : result_out = {1'b1,12'd24  };
    1029 : result_out = {1'b1,12'd30  };
    1030 : result_out = {1'b1,12'd37  };
    1031 : result_out = {1'b1,12'd43  }; 
    1032 : result_out = {1'b1,12'd49  }; 
    1033 : result_out = {1'b1,12'd56  }; 
    1034 : result_out = {1'b1,12'd62  }; 
    1035 : result_out = {1'b1,12'd68  }; 
    1036 : result_out = {1'b1,12'd74  }; 
    1037 : result_out = {1'b1,12'd81  }; 
    1038 : result_out = {1'b1,12'd87  }; 
    1039 : result_out = {1'b1,12'd93  }; 
    1040 : result_out = {1'b1,12'd100 }; 
    1041 : result_out = {1'b1,12'd106 }; 
    1042 : result_out = {1'b1,12'd112 }; 
    1043 : result_out = {1'b1,12'd118 }; 
    1044 : result_out = {1'b1,12'd125 }; 
    1045 : result_out = {1'b1,12'd131 }; 
    1046 : result_out = {1'b1,12'd137 }; 
    1047 : result_out = {1'b1,12'd143 }; 
    1048 : result_out = {1'b1,12'd150 }; 
    1049 : result_out = {1'b1,12'd156 }; 
    1050 : result_out = {1'b1,12'd162 }; 
    1051 : result_out = {1'b1,12'd169 }; 
    1052 : result_out = {1'b1,12'd175 }; 
    1053 : result_out = {1'b1,12'd181 }; 
    1054 : result_out = {1'b1,12'd187 }; 
    1055 : result_out = {1'b1,12'd194 }; 
    1056 : result_out = {1'b1,12'd200 }; 
    1057 : result_out = {1'b1,12'd206 }; 
    1058 : result_out = {1'b1,12'd213 }; 
    1059 : result_out = {1'b1,12'd219 }; 
    1060 : result_out = {1'b1,12'd225 }; 
    1061 : result_out = {1'b1,12'd231 }; 
    1062 : result_out = {1'b1,12'd238 }; 
    1063 : result_out = {1'b1,12'd244 }; 
    1064 : result_out = {1'b1,12'd250 }; 
    1065 : result_out = {1'b1,12'd256 }; 
    1066 : result_out = {1'b1,12'd263 }; 
    1067 : result_out = {1'b1,12'd269 }; 
    1068 : result_out = {1'b1,12'd275 }; 
    1069 : result_out = {1'b1,12'd282 }; 
    1070 : result_out = {1'b1,12'd288 }; 
    1071 : result_out = {1'b1,12'd294 }; 
    1072 : result_out = {1'b1,12'd300 }; 
    1073 : result_out = {1'b1,12'd307 }; 
    1074 : result_out = {1'b1,12'd313 }; 
    1075 : result_out = {1'b1,12'd319 }; 
    1076 : result_out = {1'b1,12'd325 }; 
    1077 : result_out = {1'b1,12'd332 }; 
    1078 : result_out = {1'b1,12'd338 }; 
    1079 : result_out = {1'b1,12'd344 }; 
    1080 : result_out = {1'b1,12'd350 }; 
    1081 : result_out = {1'b1,12'd357 }; 
    1082 : result_out = {1'b1,12'd363 }; 
    1083 : result_out = {1'b1,12'd369 }; 
    1084 : result_out = {1'b1,12'd375 }; 
    1085 : result_out = {1'b1,12'd382 }; 
    1086 : result_out = {1'b1,12'd388 }; 
    1087 : result_out = {1'b1,12'd394 }; 
    1088 : result_out = {1'b1,12'd400 };  
    1089 : result_out = {1'b1,12'd407 };  
    1090 : result_out = {1'b1,12'd413 };  
    1091 : result_out = {1'b1,12'd419 };  
    1092 : result_out = {1'b1,12'd425 };  
    1093 : result_out = {1'b1,12'd432 };  
    1094 : result_out = {1'b1,12'd438 };  
    1095 : result_out = {1'b1,12'd444 };  
    1096 : result_out = {1'b1,12'd450 };  
    1097 : result_out = {1'b1,12'd457 };  
    1098 : result_out = {1'b1,12'd463 };  
    1099 : result_out = {1'b1,12'd469 };  
    1100 : result_out = {1'b1,12'd475 };  
    1101 : result_out = {1'b1,12'd482 };  
    1102 : result_out = {1'b1,12'd488 };  
    1103 : result_out = {1'b1,12'd494 };  
    1104 : result_out = {1'b1,12'd500 };  
    1105 : result_out = {1'b1,12'd507 };  
    1106 : result_out = {1'b1,12'd513 };  
    1107 : result_out = {1'b1,12'd519 };  
    1108 : result_out = {1'b1,12'd525 };  
    1109 : result_out = {1'b1,12'd532 };  
    1110 : result_out = {1'b1,12'd538 };  
    1111 : result_out = {1'b1,12'd544 };  
    1112 : result_out = {1'b1,12'd550 };  
    1113 : result_out = {1'b1,12'd556 };  
    1114 : result_out = {1'b1,12'd563 };  
    1115 : result_out = {1'b1,12'd569 };  
    1116 : result_out = {1'b1,12'd575 };  
    1117 : result_out = {1'b1,12'd581 };  
    1118 : result_out = {1'b1,12'd588 };  
    1119 : result_out = {1'b1,12'd594 };  
    1120 : result_out = {1'b1,12'd600 };  
    1121 : result_out = {1'b1,12'd606 };  
    1122 : result_out = {1'b1,12'd612 };  
    1123 : result_out = {1'b1,12'd619 };  
    1124 : result_out = {1'b1,12'd625 };  
    1125 : result_out = {1'b1,12'd631 };  
    1126 : result_out = {1'b1,12'd637 };  
    1127 : result_out = {1'b1,12'd643 };  
    1128 : result_out = {1'b1,12'd650 };  
    1129 : result_out = {1'b1,12'd656 };  
    1130 : result_out = {1'b1,12'd662 };  
    1131 : result_out = {1'b1,12'd668 };  
    1132 : result_out = {1'b1,12'd674 };  
    1133 : result_out = {1'b1,12'd681 };  
    1134 : result_out = {1'b1,12'd687 };  
    1135 : result_out = {1'b1,12'd693 };  
    1136 : result_out = {1'b1,12'd699 };  
    1137 : result_out = {1'b1,12'd705 };  
    1138 : result_out = {1'b1,12'd712 };  
    1139 : result_out = {1'b1,12'd718 };  
    1140 : result_out = {1'b1,12'd724 };  
    1141 : result_out = {1'b1,12'd730 };  
    1142 : result_out = {1'b1,12'd736 };  
    1143 : result_out = {1'b1,12'd743 };  
    1144 : result_out = {1'b1,12'd749 };  
    1145 : result_out = {1'b1,12'd755 };  
    1146 : result_out = {1'b1,12'd761 };  
    1147 : result_out = {1'b1,12'd767 };  
    1148 : result_out = {1'b1,12'd773 };  
    1149 : result_out = {1'b1,12'd780 };  
    1150 : result_out = {1'b1,12'd786 };  
    1151 : result_out = {1'b1,12'd792 };  
    1152 : result_out = {1'b1,12'd798 };  
    1153 : result_out = {1'b1,12'd804 };  
    1154 : result_out = {1'b1,12'd810 };  
    1155 : result_out = {1'b1,12'd817 };  
    1156 : result_out = {1'b1,12'd823 };  
    1157 : result_out = {1'b1,12'd829 };  
    1158 : result_out = {1'b1,12'd835 };  
    1159 : result_out = {1'b1,12'd841 };  
    1160 : result_out = {1'b1,12'd847 };  
    1161 : result_out = {1'b1,12'd853 };  
    1162 : result_out = {1'b1,12'd860 };  
    1163 : result_out = {1'b1,12'd866 };  
    1164 : result_out = {1'b1,12'd872 };  
    1165 : result_out = {1'b1,12'd878 };  
    1166 : result_out = {1'b1,12'd884 };  
    1167 : result_out = {1'b1,12'd890 };  
    1168 : result_out = {1'b1,12'd896 };  
    1169 : result_out = {1'b1,12'd903 };  
    1170 : result_out = {1'b1,12'd909 };  
    1171 : result_out = {1'b1,12'd915 };  
    1172 : result_out = {1'b1,12'd921 };  
    1173 : result_out = {1'b1,12'd927 };  
    1174 : result_out = {1'b1,12'd933 };  
    1175 : result_out = {1'b1,12'd939 };  
    1176 : result_out = {1'b1,12'd945 };  
    1177 : result_out = {1'b1,12'd952 };  
    1178 : result_out = {1'b1,12'd958 };  
    1179 : result_out = {1'b1,12'd964 };  
    1180 : result_out = {1'b1,12'd970 };  
    1181 : result_out = {1'b1,12'd976 };  
    1182 : result_out = {1'b1,12'd982 };  
    1183 : result_out = {1'b1,12'd988 };  
    1184 : result_out = {1'b1,12'd994 };  
    1185 : result_out = {1'b1,12'd1000};  
    1186 : result_out = {1'b1,12'd1006};  
    1187 : result_out = {1'b1,12'd1013};  
    1188 : result_out = {1'b1,12'd1019};  
    1189 : result_out = {1'b1,12'd1025};  
    1190 : result_out = {1'b1,12'd1031};  
    1191 : result_out = {1'b1,12'd1037};  
    1192 : result_out = {1'b1,12'd1043};  
    1193 : result_out = {1'b1,12'd1049};  
    1194 : result_out = {1'b1,12'd1055};  
    1195 : result_out = {1'b1,12'd1061};  
    1196 : result_out = {1'b1,12'd1067};  
    1197 : result_out = {1'b1,12'd1073};  
    1198 : result_out = {1'b1,12'd1079};  
    1199 : result_out = {1'b1,12'd1085};  
    1200 : result_out = {1'b1,12'd1091};  
    1201 : result_out = {1'b1,12'd1098};  
    1202 : result_out = {1'b1,12'd1104};  
    1203 : result_out = {1'b1,12'd1110};  
    1204 : result_out = {1'b1,12'd1116};  
    1205 : result_out = {1'b1,12'd1122};  
    1206 : result_out = {1'b1,12'd1128};  
    1207 : result_out = {1'b1,12'd1134};  
    1208 : result_out = {1'b1,12'd1140};  
    1209 : result_out = {1'b1,12'd1146};  
    1210 : result_out = {1'b1,12'd1152};  
    1211 : result_out = {1'b1,12'd1158};  
    1212 : result_out = {1'b1,12'd1164};  
    1213 : result_out = {1'b1,12'd1170};  
    1214 : result_out = {1'b1,12'd1176};  
    1215 : result_out = {1'b1,12'd1182};  
    1216 : result_out = {1'b1,12'd1188};  
    1217 : result_out = {1'b1,12'd1194};  
    1218 : result_out = {1'b1,12'd1200};  
    1219 : result_out = {1'b1,12'd1206};  
    1220 : result_out = {1'b1,12'd1212};  
    1221 : result_out = {1'b1,12'd1218};  
    1222 : result_out = {1'b1,12'd1224};  
    1223 : result_out = {1'b1,12'd1230};  
    1224 : result_out = {1'b1,12'd1236};  
    1225 : result_out = {1'b1,12'd1242};  
    1226 : result_out = {1'b1,12'd1248};  
    1227 : result_out = {1'b1,12'd1254};  
    1228 : result_out = {1'b1,12'd1260};  
    1229 : result_out = {1'b1,12'd1266};  
    1230 : result_out = {1'b1,12'd1272};  
    1231 : result_out = {1'b1,12'd1278};  
    1232 : result_out = {1'b1,12'd1284};  
    1233 : result_out = {1'b1,12'd1290};  
    1234 : result_out = {1'b1,12'd1296};  
    1235 : result_out = {1'b1,12'd1302};  
    1236 : result_out = {1'b1,12'd1308};  
    1237 : result_out = {1'b1,12'd1314};  
    1238 : result_out = {1'b1,12'd1320};  
    1239 : result_out = {1'b1,12'd1326};  
    1240 : result_out = {1'b1,12'd1331};  
    1241 : result_out = {1'b1,12'd1337};  
    1242 : result_out = {1'b1,12'd1343};  
    1243 : result_out = {1'b1,12'd1349};  
    1244 : result_out = {1'b1,12'd1355};  
    1245 : result_out = {1'b1,12'd1361};  
    1246 : result_out = {1'b1,12'd1367};  
    1247 : result_out = {1'b1,12'd1373};  
    1248 : result_out = {1'b1,12'd1379};  
    1249 : result_out = {1'b1,12'd1385};  
    1250 : result_out = {1'b1,12'd1391};  
    1251 : result_out = {1'b1,12'd1397};  
    1252 : result_out = {1'b1,12'd1403};  
    1253 : result_out = {1'b1,12'd1408};  
    1254 : result_out = {1'b1,12'd1414};  
    1255 : result_out = {1'b1,12'd1420};  
    1256 : result_out = {1'b1,12'd1426};  
    1257 : result_out = {1'b1,12'd1432};  
    1258 : result_out = {1'b1,12'd1438};  
    1259 : result_out = {1'b1,12'd1444};  
    1260 : result_out = {1'b1,12'd1450};  
    1261 : result_out = {1'b1,12'd1456};  
    1262 : result_out = {1'b1,12'd1461};  
    1263 : result_out = {1'b1,12'd1467};  
    1264 : result_out = {1'b1,12'd1473};  
    1265 : result_out = {1'b1,12'd1479};  
    1266 : result_out = {1'b1,12'd1485};  
    1267 : result_out = {1'b1,12'd1491};  
    1268 : result_out = {1'b1,12'd1497};  
    1269 : result_out = {1'b1,12'd1502};  
    1270 : result_out = {1'b1,12'd1508};  
    1271 : result_out = {1'b1,12'd1514};  
    1272 : result_out = {1'b1,12'd1520};  
    1273 : result_out = {1'b1,12'd1526};  
    1274 : result_out = {1'b1,12'd1532};  
    1275 : result_out = {1'b1,12'd1537};  
    1276 : result_out = {1'b1,12'd1543};  
    1277 : result_out = {1'b1,12'd1549};  
    1278 : result_out = {1'b1,12'd1555};  
    1279 : result_out = {1'b1,12'd1561};  
    1280 : result_out = {1'b1,12'd1566};  
    1281 : result_out = {1'b1,12'd1572};  
    1282 : result_out = {1'b1,12'd1578};  
    1283 : result_out = {1'b1,12'd1584};  
    1284 : result_out = {1'b1,12'd1590};  
    1285 : result_out = {1'b1,12'd1595};  
    1286 : result_out = {1'b1,12'd1601};  
    1287 : result_out = {1'b1,12'd1607};  
    1288 : result_out = {1'b1,12'd1613};  
    1289 : result_out = {1'b1,12'd1619};  
    1290 : result_out = {1'b1,12'd1624};  
    1291 : result_out = {1'b1,12'd1630};  
    1292 : result_out = {1'b1,12'd1636};  
    1293 : result_out = {1'b1,12'd1642};  
    1294 : result_out = {1'b1,12'd1647};  
    1295 : result_out = {1'b1,12'd1653};  
    1296 : result_out = {1'b1,12'd1659};  
    1297 : result_out = {1'b1,12'd1665};  
    1298 : result_out = {1'b1,12'd1670};  
    1299 : result_out = {1'b1,12'd1676};  
    1300 : result_out = {1'b1,12'd1682};  
    1301 : result_out = {1'b1,12'd1688};  
    1302 : result_out = {1'b1,12'd1693};  
    1303 : result_out = {1'b1,12'd1699};  
    1304 : result_out = {1'b1,12'd1705};  
    1305 : result_out = {1'b1,12'd1710};  
    1306 : result_out = {1'b1,12'd1716};  
    1307 : result_out = {1'b1,12'd1722};  
    1308 : result_out = {1'b1,12'd1728};  
    1309 : result_out = {1'b1,12'd1733};  
    1310 : result_out = {1'b1,12'd1739};  
    1311 : result_out = {1'b1,12'd1745};  
    1312 : result_out = {1'b1,12'd1750};  
    1313 : result_out = {1'b1,12'd1756};  
    1314 : result_out = {1'b1,12'd1762};  
    1315 : result_out = {1'b1,12'd1767};  
    1316 : result_out = {1'b1,12'd1773};  
    1317 : result_out = {1'b1,12'd1779};  
    1318 : result_out = {1'b1,12'd1784};  
    1319 : result_out = {1'b1,12'd1790};  
    1320 : result_out = {1'b1,12'd1796};  
    1321 : result_out = {1'b1,12'd1801};  
    1322 : result_out = {1'b1,12'd1807};  
    1323 : result_out = {1'b1,12'd1812};  
    1324 : result_out = {1'b1,12'd1818};  
    1325 : result_out = {1'b1,12'd1824};  
    1326 : result_out = {1'b1,12'd1829};  
    1327 : result_out = {1'b1,12'd1835};  
    1328 : result_out = {1'b1,12'd1841};  
    1329 : result_out = {1'b1,12'd1846};  
    1330 : result_out = {1'b1,12'd1852};  
    1331 : result_out = {1'b1,12'd1857};  
    1332 : result_out = {1'b1,12'd1863};  
    1333 : result_out = {1'b1,12'd1869};  
    1334 : result_out = {1'b1,12'd1874};  
    1335 : result_out = {1'b1,12'd1880};  
    1336 : result_out = {1'b1,12'd1885};  
    1337 : result_out = {1'b1,12'd1891};  
    1338 : result_out = {1'b1,12'd1897};  
    1339 : result_out = {1'b1,12'd1902};  
    1340 : result_out = {1'b1,12'd1908};  
    1341 : result_out = {1'b1,12'd1913};  
    1342 : result_out = {1'b1,12'd1919};  
    1343 : result_out = {1'b1,12'd1924};  
    1344 : result_out = {1'b1,12'd1930};  
    1345 : result_out = {1'b1,12'd1935};  
    1346 : result_out = {1'b1,12'd1941};  
    1347 : result_out = {1'b1,12'd1946};  
    1348 : result_out = {1'b1,12'd1952};  
    1349 : result_out = {1'b1,12'd1957};  
    1350 : result_out = {1'b1,12'd1963};  
    1351 : result_out = {1'b1,12'd1969};  
    1352 : result_out = {1'b1,12'd1974};  
    1353 : result_out = {1'b1,12'd1980};  
    1354 : result_out = {1'b1,12'd1985};  
    1355 : result_out = {1'b1,12'd1991};  
    1356 : result_out = {1'b1,12'd1996};  
    1357 : result_out = {1'b1,12'd2001};  
    1358 : result_out = {1'b1,12'd2007};  
    1359 : result_out = {1'b1,12'd2012};  
    1360 : result_out = {1'b1,12'd2018};  
    1361 : result_out = {1'b1,12'd2023};  
    1362 : result_out = {1'b1,12'd2029};  
    1363 : result_out = {1'b1,12'd2034};  
    1364 : result_out = {1'b1,12'd2040};  
    1365 : result_out = {1'b1,12'd2045};  
    1366 : result_out = {1'b1,12'd2051};  
    1367 : result_out = {1'b1,12'd2056};  
    1368 : result_out = {1'b1,12'd2061};  
    1369 : result_out = {1'b1,12'd2067};  
    1370 : result_out = {1'b1,12'd2072};  
    1371 : result_out = {1'b1,12'd2078};  
    1372 : result_out = {1'b1,12'd2083};  
    1373 : result_out = {1'b1,12'd2089};  
    1374 : result_out = {1'b1,12'd2094};  
    1375 : result_out = {1'b1,12'd2099};  
    1376 : result_out = {1'b1,12'd2105};  
    1377 : result_out = {1'b1,12'd2110};  
    1378 : result_out = {1'b1,12'd2116};  
    1379 : result_out = {1'b1,12'd2121};  
    1380 : result_out = {1'b1,12'd2126};  
    1381 : result_out = {1'b1,12'd2132};  
    1382 : result_out = {1'b1,12'd2137};  
    1383 : result_out = {1'b1,12'd2142};  
    1384 : result_out = {1'b1,12'd2148};  
    1385 : result_out = {1'b1,12'd2153};  
    1386 : result_out = {1'b1,12'd2158};  
    1387 : result_out = {1'b1,12'd2164};  
    1388 : result_out = {1'b1,12'd2169};  
    1389 : result_out = {1'b1,12'd2174};  
    1390 : result_out = {1'b1,12'd2180};  
    1391 : result_out = {1'b1,12'd2185};  
    1392 : result_out = {1'b1,12'd2190};  
    1393 : result_out = {1'b1,12'd2196};  
    1394 : result_out = {1'b1,12'd2201};  
    1395 : result_out = {1'b1,12'd2206};  
    1396 : result_out = {1'b1,12'd2212};  
    1397 : result_out = {1'b1,12'd2217};  
    1398 : result_out = {1'b1,12'd2222};  
    1399 : result_out = {1'b1,12'd2227};  
    1400 : result_out = {1'b1,12'd2233};  
    1401 : result_out = {1'b1,12'd2238};  
    1402 : result_out = {1'b1,12'd2243};  
    1403 : result_out = {1'b1,12'd2248};  
    1404 : result_out = {1'b1,12'd2254};  
    1405 : result_out = {1'b1,12'd2259};  
    1406 : result_out = {1'b1,12'd2264};  
    1407 : result_out = {1'b1,12'd2269};  
    1408 : result_out = {1'b1,12'd2275};  
    1409 : result_out = {1'b1,12'd2280};  
    1410 : result_out = {1'b1,12'd2285};  
    1411 : result_out = {1'b1,12'd2290};  
    1412 : result_out = {1'b1,12'd2295};  
    1413 : result_out = {1'b1,12'd2301};  
    1414 : result_out = {1'b1,12'd2306};  
    1415 : result_out = {1'b1,12'd2311};  
    1416 : result_out = {1'b1,12'd2316};  
    1417 : result_out = {1'b1,12'd2321};  
    1418 : result_out = {1'b1,12'd2327};  
    1419 : result_out = {1'b1,12'd2332};  
    1420 : result_out = {1'b1,12'd2337};  
    1421 : result_out = {1'b1,12'd2342};  
    1422 : result_out = {1'b1,12'd2347};  
    1423 : result_out = {1'b1,12'd2352};  
    1424 : result_out = {1'b1,12'd2358};  
    1425 : result_out = {1'b1,12'd2363};  
    1426 : result_out = {1'b1,12'd2368};  
    1427 : result_out = {1'b1,12'd2373};  
    1428 : result_out = {1'b1,12'd2378};  
    1429 : result_out = {1'b1,12'd2383};  
    1430 : result_out = {1'b1,12'd2388};  
    1431 : result_out = {1'b1,12'd2393};  
    1432 : result_out = {1'b1,12'd2398};  
    1433 : result_out = {1'b1,12'd2404};  
    1434 : result_out = {1'b1,12'd2409};  
    1435 : result_out = {1'b1,12'd2414};  
    1436 : result_out = {1'b1,12'd2419};  
    1437 : result_out = {1'b1,12'd2424};  
    1438 : result_out = {1'b1,12'd2429};  
    1439 : result_out = {1'b1,12'd2434};  
    1440 : result_out = {1'b1,12'd2439};  
    1441 : result_out = {1'b1,12'd2444};  
    1442 : result_out = {1'b1,12'd2449};  
    1443 : result_out = {1'b1,12'd2454};  
    1444 : result_out = {1'b1,12'd2459};  
    1445 : result_out = {1'b1,12'd2464};  
    1446 : result_out = {1'b1,12'd2469};  
    1447 : result_out = {1'b1,12'd2474};  
    1448 : result_out = {1'b1,12'd2479};  
    1449 : result_out = {1'b1,12'd2484};  
    1450 : result_out = {1'b1,12'd2489};  
    1451 : result_out = {1'b1,12'd2494};  
    1452 : result_out = {1'b1,12'd2499};  
    1453 : result_out = {1'b1,12'd2504};  
    1454 : result_out = {1'b1,12'd2509};  
    1455 : result_out = {1'b1,12'd2514};  
    1456 : result_out = {1'b1,12'd2519};  
    1457 : result_out = {1'b1,12'd2524};  
    1458 : result_out = {1'b1,12'd2529};  
    1459 : result_out = {1'b1,12'd2534};  
    1460 : result_out = {1'b1,12'd2539};  
    1461 : result_out = {1'b1,12'd2544};  
    1462 : result_out = {1'b1,12'd2549};  
    1463 : result_out = {1'b1,12'd2554};  
    1464 : result_out = {1'b1,12'd2558};  
    1465 : result_out = {1'b1,12'd2563};  
    1466 : result_out = {1'b1,12'd2568};  
    1467 : result_out = {1'b1,12'd2573};  
    1468 : result_out = {1'b1,12'd2578};  
    1469 : result_out = {1'b1,12'd2583};  
    1470 : result_out = {1'b1,12'd2588};  
    1471 : result_out = {1'b1,12'd2593};  
    1472 : result_out = {1'b1,12'd2597};  
    1473 : result_out = {1'b1,12'd2602};  
    1474 : result_out = {1'b1,12'd2607};  
    1475 : result_out = {1'b1,12'd2612};  
    1476 : result_out = {1'b1,12'd2617};  
    1477 : result_out = {1'b1,12'd2622};  
    1478 : result_out = {1'b1,12'd2627};  
    1479 : result_out = {1'b1,12'd2631};  
    1480 : result_out = {1'b1,12'd2636};  
    1481 : result_out = {1'b1,12'd2641};  
    1482 : result_out = {1'b1,12'd2646};  
    1483 : result_out = {1'b1,12'd2651};  
    1484 : result_out = {1'b1,12'd2655};  
    1485 : result_out = {1'b1,12'd2660};  
    1486 : result_out = {1'b1,12'd2665};  
    1487 : result_out = {1'b1,12'd2670};  
    1488 : result_out = {1'b1,12'd2674};  
    1489 : result_out = {1'b1,12'd2679};  
    1490 : result_out = {1'b1,12'd2684};  
    1491 : result_out = {1'b1,12'd2689};  
    1492 : result_out = {1'b1,12'd2693};  
    1493 : result_out = {1'b1,12'd2698};  
    1494 : result_out = {1'b1,12'd2703};  
    1495 : result_out = {1'b1,12'd2708};  
    1496 : result_out = {1'b1,12'd2712};  
    1497 : result_out = {1'b1,12'd2717};  
    1498 : result_out = {1'b1,12'd2722};  
    1499 : result_out = {1'b1,12'd2726};  
    1500 : result_out = {1'b1,12'd2731};  
    1501 : result_out = {1'b1,12'd2736};  
    1502 : result_out = {1'b1,12'd2740};  
    1503 : result_out = {1'b1,12'd2745};  
    1504 : result_out = {1'b1,12'd2750};  
    1505 : result_out = {1'b1,12'd2754};  
    1506 : result_out = {1'b1,12'd2759};  
    1507 : result_out = {1'b1,12'd2764};  
    1508 : result_out = {1'b1,12'd2768};  
    1509 : result_out = {1'b1,12'd2773};  
    1510 : result_out = {1'b1,12'd2778};  
    1511 : result_out = {1'b1,12'd2782};  
    1512 : result_out = {1'b1,12'd2787};  
    1513 : result_out = {1'b1,12'd2791};  
    1514 : result_out = {1'b1,12'd2796};  
    1515 : result_out = {1'b1,12'd2801};  
    1516 : result_out = {1'b1,12'd2805};  
    1517 : result_out = {1'b1,12'd2810};  
    1518 : result_out = {1'b1,12'd2814};  
    1519 : result_out = {1'b1,12'd2819};  
    1520 : result_out = {1'b1,12'd2823};  
    1521 : result_out = {1'b1,12'd2828};  
    1522 : result_out = {1'b1,12'd2832};  
    1523 : result_out = {1'b1,12'd2837};  
    1524 : result_out = {1'b1,12'd2842};  
    1525 : result_out = {1'b1,12'd2846};  
    1526 : result_out = {1'b1,12'd2851};  
    1527 : result_out = {1'b1,12'd2855};  
    1528 : result_out = {1'b1,12'd2860};  
    1529 : result_out = {1'b1,12'd2864};  
    1530 : result_out = {1'b1,12'd2869};  
    1531 : result_out = {1'b1,12'd2873};  
    1532 : result_out = {1'b1,12'd2877};  
    1533 : result_out = {1'b1,12'd2882};  
    1534 : result_out = {1'b1,12'd2886};  
    1535 : result_out = {1'b1,12'd2891};  
    1536 : result_out = {1'b1,12'd2895};  
    1537 : result_out = {1'b1,12'd2900};  
    1538 : result_out = {1'b1,12'd2904};  
    1539 : result_out = {1'b1,12'd2909};  
    1540 : result_out = {1'b1,12'd2913};  
    1541 : result_out = {1'b1,12'd2917};  
    1542 : result_out = {1'b1,12'd2922};  
    1543 : result_out = {1'b1,12'd2926};  
    1544 : result_out = {1'b1,12'd2931};  
    1545 : result_out = {1'b1,12'd2935};  
    1546 : result_out = {1'b1,12'd2939};  
    1547 : result_out = {1'b1,12'd2944};  
    1548 : result_out = {1'b1,12'd2948};  
    1549 : result_out = {1'b1,12'd2952};  
    1550 : result_out = {1'b1,12'd2957};  
    1551 : result_out = {1'b1,12'd2961};  
    1552 : result_out = {1'b1,12'd2966};  
    1553 : result_out = {1'b1,12'd2970};  
    1554 : result_out = {1'b1,12'd2974};  
    1555 : result_out = {1'b1,12'd2978};  
    1556 : result_out = {1'b1,12'd2983};  
    1557 : result_out = {1'b1,12'd2987};  
    1558 : result_out = {1'b1,12'd2991};  
    1559 : result_out = {1'b1,12'd2996};  
    1560 : result_out = {1'b1,12'd3000};  
    1561 : result_out = {1'b1,12'd3004};  
    1562 : result_out = {1'b1,12'd3008};  
    1563 : result_out = {1'b1,12'd3013};  
    1564 : result_out = {1'b1,12'd3017};  
    1565 : result_out = {1'b1,12'd3021};  
    1566 : result_out = {1'b1,12'd3025};  
    1567 : result_out = {1'b1,12'd3030};  
    1568 : result_out = {1'b1,12'd3034};  
    1569 : result_out = {1'b1,12'd3038};  
    1570 : result_out = {1'b1,12'd3042};  
    1571 : result_out = {1'b1,12'd3047};  
    1572 : result_out = {1'b1,12'd3051};  
    1573 : result_out = {1'b1,12'd3055};  
    1574 : result_out = {1'b1,12'd3059};  
    1575 : result_out = {1'b1,12'd3063};  
    1576 : result_out = {1'b1,12'd3067};  
    1577 : result_out = {1'b1,12'd3072};  
    1578 : result_out = {1'b1,12'd3076};  
    1579 : result_out = {1'b1,12'd3080};  
    1580 : result_out = {1'b1,12'd3084};  
    1581 : result_out = {1'b1,12'd3088};  
    1582 : result_out = {1'b1,12'd3092};  
    1583 : result_out = {1'b1,12'd3096};  
    1584 : result_out = {1'b1,12'd3101};  
    1585 : result_out = {1'b1,12'd3105};  
    1586 : result_out = {1'b1,12'd3109};  
    1587 : result_out = {1'b1,12'd3113};  
    1588 : result_out = {1'b1,12'd3117};  
    1589 : result_out = {1'b1,12'd3121};  
    1590 : result_out = {1'b1,12'd3125};  
    1591 : result_out = {1'b1,12'd3129};  
    1592 : result_out = {1'b1,12'd3133};  
    1593 : result_out = {1'b1,12'd3137};  
    1594 : result_out = {1'b1,12'd3141};  
    1595 : result_out = {1'b1,12'd3145};  
    1596 : result_out = {1'b1,12'd3149};  
    1597 : result_out = {1'b1,12'd3153};  
    1598 : result_out = {1'b1,12'd3157};  
    1599 : result_out = {1'b1,12'd3161};  
    1600 : result_out = {1'b1,12'd3165};  
    1601 : result_out = {1'b1,12'd3169};  
    1602 : result_out = {1'b1,12'd3173};  
    1603 : result_out = {1'b1,12'd3177};  
    1604 : result_out = {1'b1,12'd3181};  
    1605 : result_out = {1'b1,12'd3185};  
    1606 : result_out = {1'b1,12'd3189};  
    1607 : result_out = {1'b1,12'd3193};  
    1608 : result_out = {1'b1,12'd3197};  
    1609 : result_out = {1'b1,12'd3201};  
    1610 : result_out = {1'b1,12'd3205};  
    1611 : result_out = {1'b1,12'd3209};  
    1612 : result_out = {1'b1,12'd3213};  
    1613 : result_out = {1'b1,12'd3216};  
    1614 : result_out = {1'b1,12'd3220};  
    1615 : result_out = {1'b1,12'd3224};  
    1616 : result_out = {1'b1,12'd3228};  
    1617 : result_out = {1'b1,12'd3232};  
    1618 : result_out = {1'b1,12'd3236};  
    1619 : result_out = {1'b1,12'd3240};  
    1620 : result_out = {1'b1,12'd3243};  
    1621 : result_out = {1'b1,12'd3247};  
    1622 : result_out = {1'b1,12'd3251};  
    1623 : result_out = {1'b1,12'd3255};  
    1624 : result_out = {1'b1,12'd3259};  
    1625 : result_out = {1'b1,12'd3263};  
    1626 : result_out = {1'b1,12'd3266};  
    1627 : result_out = {1'b1,12'd3270};  
    1628 : result_out = {1'b1,12'd3274};  
    1629 : result_out = {1'b1,12'd3278};  
    1630 : result_out = {1'b1,12'd3281};  
    1631 : result_out = {1'b1,12'd3285};  
    1632 : result_out = {1'b1,12'd3289};  
    1633 : result_out = {1'b1,12'd3293};  
    1634 : result_out = {1'b1,12'd3296};  
    1635 : result_out = {1'b1,12'd3300};  
    1636 : result_out = {1'b1,12'd3304};  
    1637 : result_out = {1'b1,12'd3308};  
    1638 : result_out = {1'b1,12'd3311};  
    1639 : result_out = {1'b1,12'd3315};  
    1640 : result_out = {1'b1,12'd3319};  
    1641 : result_out = {1'b1,12'd3322};  
    1642 : result_out = {1'b1,12'd3326};  
    1643 : result_out = {1'b1,12'd3330};  
    1644 : result_out = {1'b1,12'd3333};  
    1645 : result_out = {1'b1,12'd3337};  
    1646 : result_out = {1'b1,12'd3341};  
    1647 : result_out = {1'b1,12'd3344};  
    1648 : result_out = {1'b1,12'd3348};  
    1649 : result_out = {1'b1,12'd3351};  
    1650 : result_out = {1'b1,12'd3355};  
    1651 : result_out = {1'b1,12'd3359};  
    1652 : result_out = {1'b1,12'd3362};  
    1653 : result_out = {1'b1,12'd3366};  
    1654 : result_out = {1'b1,12'd3369};  
    1655 : result_out = {1'b1,12'd3373};  
    1656 : result_out = {1'b1,12'd3377};  
    1657 : result_out = {1'b1,12'd3380};  
    1658 : result_out = {1'b1,12'd3384};  
    1659 : result_out = {1'b1,12'd3387};  
    1660 : result_out = {1'b1,12'd3391};  
    1661 : result_out = {1'b1,12'd3394};  
    1662 : result_out = {1'b1,12'd3398};  
    1663 : result_out = {1'b1,12'd3401};  
    1664 : result_out = {1'b1,12'd3405};  
    1665 : result_out = {1'b1,12'd3408};  
    1666 : result_out = {1'b1,12'd3412};  
    1667 : result_out = {1'b1,12'd3415};  
    1668 : result_out = {1'b1,12'd3419};  
    1669 : result_out = {1'b1,12'd3422};  
    1670 : result_out = {1'b1,12'd3425};  
    1671 : result_out = {1'b1,12'd3429};  
    1672 : result_out = {1'b1,12'd3432};  
    1673 : result_out = {1'b1,12'd3436};  
    1674 : result_out = {1'b1,12'd3439};  
    1675 : result_out = {1'b1,12'd3443};  
    1676 : result_out = {1'b1,12'd3446};  
    1677 : result_out = {1'b1,12'd3449};  
    1678 : result_out = {1'b1,12'd3453};  
    1679 : result_out = {1'b1,12'd3456};  
    1680 : result_out = {1'b1,12'd3460};  
    1681 : result_out = {1'b1,12'd3463};  
    1682 : result_out = {1'b1,12'd3466};  
    1683 : result_out = {1'b1,12'd3470};  
    1684 : result_out = {1'b1,12'd3473};  
    1685 : result_out = {1'b1,12'd3476};  
    1686 : result_out = {1'b1,12'd3480};  
    1687 : result_out = {1'b1,12'd3483};  
    1688 : result_out = {1'b1,12'd3486};  
    1689 : result_out = {1'b1,12'd3489};  
    1690 : result_out = {1'b1,12'd3493};  
    1691 : result_out = {1'b1,12'd3496};  
    1692 : result_out = {1'b1,12'd3499};  
    1693 : result_out = {1'b1,12'd3503};  
    1694 : result_out = {1'b1,12'd3506};  
    1695 : result_out = {1'b1,12'd3509};  
    1696 : result_out = {1'b1,12'd3512};  
    1697 : result_out = {1'b1,12'd3515};  
    1698 : result_out = {1'b1,12'd3519};  
    1699 : result_out = {1'b1,12'd3522};  
    1700 : result_out = {1'b1,12'd3525};  
    1701 : result_out = {1'b1,12'd3528};  
    1702 : result_out = {1'b1,12'd3531};  
    1703 : result_out = {1'b1,12'd3535};  
    1704 : result_out = {1'b1,12'd3538};  
    1705 : result_out = {1'b1,12'd3541};  
    1706 : result_out = {1'b1,12'd3544};  
    1707 : result_out = {1'b1,12'd3547};  
    1708 : result_out = {1'b1,12'd3550};  
    1709 : result_out = {1'b1,12'd3554};  
    1710 : result_out = {1'b1,12'd3557};  
    1711 : result_out = {1'b1,12'd3560};  
    1712 : result_out = {1'b1,12'd3563};  
    1713 : result_out = {1'b1,12'd3566};  
    1714 : result_out = {1'b1,12'd3569};  
    1715 : result_out = {1'b1,12'd3572};  
    1716 : result_out = {1'b1,12'd3575};  
    1717 : result_out = {1'b1,12'd3578};  
    1718 : result_out = {1'b1,12'd3581};  
    1719 : result_out = {1'b1,12'd3584};  
    1720 : result_out = {1'b1,12'd3587};  
    1721 : result_out = {1'b1,12'd3590};  
    1722 : result_out = {1'b1,12'd3593};  
    1723 : result_out = {1'b1,12'd3596};  
    1724 : result_out = {1'b1,12'd3599};  
    1725 : result_out = {1'b1,12'd3602};  
    1726 : result_out = {1'b1,12'd3605};  
    1727 : result_out = {1'b1,12'd3608};  
    1728 : result_out = {1'b1,12'd3611};  
    1729 : result_out = {1'b1,12'd3614};  
    1730 : result_out = {1'b1,12'd3617};  
    1731 : result_out = {1'b1,12'd3620};  
    1732 : result_out = {1'b1,12'd3623};  
    1733 : result_out = {1'b1,12'd3626};  
    1734 : result_out = {1'b1,12'd3629};  
    1735 : result_out = {1'b1,12'd3632};  
    1736 : result_out = {1'b1,12'd3635};  
    1737 : result_out = {1'b1,12'd3638};  
    1738 : result_out = {1'b1,12'd3641};  
    1739 : result_out = {1'b1,12'd3643};  
    1740 : result_out = {1'b1,12'd3646};  
    1741 : result_out = {1'b1,12'd3649};  
    1742 : result_out = {1'b1,12'd3652};  
    1743 : result_out = {1'b1,12'd3655};  
    1744 : result_out = {1'b1,12'd3658};  
    1745 : result_out = {1'b1,12'd3660};  
    1746 : result_out = {1'b1,12'd3663};  
    1747 : result_out = {1'b1,12'd3666};  
    1748 : result_out = {1'b1,12'd3669};  
    1749 : result_out = {1'b1,12'd3672};  
    1750 : result_out = {1'b1,12'd3674};  
    1751 : result_out = {1'b1,12'd3677};  
    1752 : result_out = {1'b1,12'd3680};  
    1753 : result_out = {1'b1,12'd3683};  
    1754 : result_out = {1'b1,12'd3685};  
    1755 : result_out = {1'b1,12'd3688};  
    1756 : result_out = {1'b1,12'd3691};  
    1757 : result_out = {1'b1,12'd3694};  
    1758 : result_out = {1'b1,12'd3696};  
    1759 : result_out = {1'b1,12'd3699};  
    1760 : result_out = {1'b1,12'd3702};  
    1761 : result_out = {1'b1,12'd3704};  
    1762 : result_out = {1'b1,12'd3707};  
    1763 : result_out = {1'b1,12'd3710};  
    1764 : result_out = {1'b1,12'd3712};  
    1765 : result_out = {1'b1,12'd3715};  
    1766 : result_out = {1'b1,12'd3718};  
    1767 : result_out = {1'b1,12'd3720};  
    1768 : result_out = {1'b1,12'd3723};  
    1769 : result_out = {1'b1,12'd3726};  
    1770 : result_out = {1'b1,12'd3728};  
    1771 : result_out = {1'b1,12'd3731};  
    1772 : result_out = {1'b1,12'd3733};  
    1773 : result_out = {1'b1,12'd3736};  
    1774 : result_out = {1'b1,12'd3738};  
    1775 : result_out = {1'b1,12'd3741};  
    1776 : result_out = {1'b1,12'd3744};  
    1777 : result_out = {1'b1,12'd3746};  
    1778 : result_out = {1'b1,12'd3749};  
    1779 : result_out = {1'b1,12'd3751};  
    1780 : result_out = {1'b1,12'd3754};  
    1781 : result_out = {1'b1,12'd3756};  
    1782 : result_out = {1'b1,12'd3759};  
    1783 : result_out = {1'b1,12'd3761};  
    1784 : result_out = {1'b1,12'd3764};  
    1785 : result_out = {1'b1,12'd3766};  
    1786 : result_out = {1'b1,12'd3769};  
    1787 : result_out = {1'b1,12'd3771};  
    1788 : result_out = {1'b1,12'd3774};  
    1789 : result_out = {1'b1,12'd3776};  
    1790 : result_out = {1'b1,12'd3778};  
    1791 : result_out = {1'b1,12'd3781};  
    1792 : result_out = {1'b1,12'd3783};  
    1793 : result_out = {1'b1,12'd3786};  
    1794 : result_out = {1'b1,12'd3788};  
    1795 : result_out = {1'b1,12'd3790};  
    1796 : result_out = {1'b1,12'd3793};  
    1797 : result_out = {1'b1,12'd3795};  
    1798 : result_out = {1'b1,12'd3797};  
    1799 : result_out = {1'b1,12'd3800};  
    1800 : result_out = {1'b1,12'd3802};  
    1801 : result_out = {1'b1,12'd3804};  
    1802 : result_out = {1'b1,12'd3807};  
    1803 : result_out = {1'b1,12'd3809};  
    1804 : result_out = {1'b1,12'd3811};  
    1805 : result_out = {1'b1,12'd3814};  
    1806 : result_out = {1'b1,12'd3816};  
    1807 : result_out = {1'b1,12'd3818};  
    1808 : result_out = {1'b1,12'd3821};  
    1809 : result_out = {1'b1,12'd3823};  
    1810 : result_out = {1'b1,12'd3825};  
    1811 : result_out = {1'b1,12'd3827};  
    1812 : result_out = {1'b1,12'd3830};  
    1813 : result_out = {1'b1,12'd3832};  
    1814 : result_out = {1'b1,12'd3834};  
    1815 : result_out = {1'b1,12'd3836};  
    1816 : result_out = {1'b1,12'd3838};  
    1817 : result_out = {1'b1,12'd3841};  
    1818 : result_out = {1'b1,12'd3843};  
    1819 : result_out = {1'b1,12'd3845};  
    1820 : result_out = {1'b1,12'd3847};  
    1821 : result_out = {1'b1,12'd3849};  
    1822 : result_out = {1'b1,12'd3851};  
    1823 : result_out = {1'b1,12'd3853};  
    1824 : result_out = {1'b1,12'd3856};  
    1825 : result_out = {1'b1,12'd3858};  
    1826 : result_out = {1'b1,12'd3860};  
    1827 : result_out = {1'b1,12'd3862};  
    1828 : result_out = {1'b1,12'd3864};  
    1829 : result_out = {1'b1,12'd3866};  
    1830 : result_out = {1'b1,12'd3868};  
    1831 : result_out = {1'b1,12'd3870};  
    1832 : result_out = {1'b1,12'd3872};  
    1833 : result_out = {1'b1,12'd3874};  
    1834 : result_out = {1'b1,12'd3876};  
    1835 : result_out = {1'b1,12'd3878};  
    1836 : result_out = {1'b1,12'd3880};  
    1837 : result_out = {1'b1,12'd3882};  
    1838 : result_out = {1'b1,12'd3884};  
    1839 : result_out = {1'b1,12'd3886};  
    1840 : result_out = {1'b1,12'd3888};  
    1841 : result_out = {1'b1,12'd3890};  
    1842 : result_out = {1'b1,12'd3892};  
    1843 : result_out = {1'b1,12'd3894};  
    1844 : result_out = {1'b1,12'd3896};  
    1845 : result_out = {1'b1,12'd3898};  
    1846 : result_out = {1'b1,12'd3900};  
    1847 : result_out = {1'b1,12'd3902};  
    1848 : result_out = {1'b1,12'd3904};  
    1849 : result_out = {1'b1,12'd3906};  
    1850 : result_out = {1'b1,12'd3908};  
    1851 : result_out = {1'b1,12'd3909};  
    1852 : result_out = {1'b1,12'd3911};  
    1853 : result_out = {1'b1,12'd3913};  
    1854 : result_out = {1'b1,12'd3915};  
    1855 : result_out = {1'b1,12'd3917};  
    1856 : result_out = {1'b1,12'd3919};  
    1857 : result_out = {1'b1,12'd3920};  
    1858 : result_out = {1'b1,12'd3922};  
    1859 : result_out = {1'b1,12'd3924};  
    1860 : result_out = {1'b1,12'd3926};  
    1861 : result_out = {1'b1,12'd3928};  
    1862 : result_out = {1'b1,12'd3929};  
    1863 : result_out = {1'b1,12'd3931};  
    1864 : result_out = {1'b1,12'd3933};  
    1865 : result_out = {1'b1,12'd3935};  
    1866 : result_out = {1'b1,12'd3936};  
    1867 : result_out = {1'b1,12'd3938};  
    1868 : result_out = {1'b1,12'd3940};  
    1869 : result_out = {1'b1,12'd3942};  
    1870 : result_out = {1'b1,12'd3943};  
    1871 : result_out = {1'b1,12'd3945};  
    1872 : result_out = {1'b1,12'd3947};  
    1873 : result_out = {1'b1,12'd3948};  
    1874 : result_out = {1'b1,12'd3950};  
    1875 : result_out = {1'b1,12'd3952};  
    1876 : result_out = {1'b1,12'd3953};  
    1877 : result_out = {1'b1,12'd3955};  
    1878 : result_out = {1'b1,12'd3957};  
    1879 : result_out = {1'b1,12'd3958};  
    1880 : result_out = {1'b1,12'd3960};  
    1881 : result_out = {1'b1,12'd3961};  
    1882 : result_out = {1'b1,12'd3963};  
    1883 : result_out = {1'b1,12'd3964};  
    1884 : result_out = {1'b1,12'd3966};  
    1885 : result_out = {1'b1,12'd3968};  
    1886 : result_out = {1'b1,12'd3969};  
    1887 : result_out = {1'b1,12'd3971};  
    1888 : result_out = {1'b1,12'd3972};  
    1889 : result_out = {1'b1,12'd3974};  
    1890 : result_out = {1'b1,12'd3975};  
    1891 : result_out = {1'b1,12'd3977};  
    1892 : result_out = {1'b1,12'd3978};  
    1893 : result_out = {1'b1,12'd3980};  
    1894 : result_out = {1'b1,12'd3981};  
    1895 : result_out = {1'b1,12'd3983};  
    1896 : result_out = {1'b1,12'd3984};  
    1897 : result_out = {1'b1,12'd3986};  
    1898 : result_out = {1'b1,12'd3987};  
    1899 : result_out = {1'b1,12'd3988};  
    1900 : result_out = {1'b1,12'd3990};  
    1901 : result_out = {1'b1,12'd3991};  
    1902 : result_out = {1'b1,12'd3993};  
    1903 : result_out = {1'b1,12'd3994};  
    1904 : result_out = {1'b1,12'd3995};  
    1905 : result_out = {1'b1,12'd3997};  
    1906 : result_out = {1'b1,12'd3998};   
    1907 : result_out = {1'b1,12'd4000};   
    1908 : result_out = {1'b1,12'd4001};   
    1909 : result_out = {1'b1,12'd4002};   
    1910 : result_out = {1'b1,12'd4004};   
    1911 : result_out = {1'b1,12'd4005};   
    1912 : result_out = {1'b1,12'd4006};   
    1913 : result_out = {1'b1,12'd4007};   
    1914 : result_out = {1'b1,12'd4009};   
    1915 : result_out = {1'b1,12'd4010};   
    1916 : result_out = {1'b1,12'd4011};   
    1917 : result_out = {1'b1,12'd4013};   
    1918 : result_out = {1'b1,12'd4014};   
    1919 : result_out = {1'b1,12'd4015};   
    1920 : result_out = {1'b1,12'd4016};   
    1921 : result_out = {1'b1,12'd4018};   
    1922 : result_out = {1'b1,12'd4019};   
    1923 : result_out = {1'b1,12'd4020};   
    1924 : result_out = {1'b1,12'd4021};   
    1925 : result_out = {1'b1,12'd4022};   
    1926 : result_out = {1'b1,12'd4023};   
    1927 : result_out = {1'b1,12'd4025};   
    1928 : result_out = {1'b1,12'd4026};   
    1929 : result_out = {1'b1,12'd4027};   
    1930 : result_out = {1'b1,12'd4028};   
    1931 : result_out = {1'b1,12'd4029};   
    1932 : result_out = {1'b1,12'd4030};   
    1933 : result_out = {1'b1,12'd4031};   
    1934 : result_out = {1'b1,12'd4033};   
    1935 : result_out = {1'b1,12'd4034};   
    1936 : result_out = {1'b1,12'd4035};   
    1937 : result_out = {1'b1,12'd4036};   
    1938 : result_out = {1'b1,12'd4037};   
    1939 : result_out = {1'b1,12'd4038};   
    1940 : result_out = {1'b1,12'd4039};   
    1941 : result_out = {1'b1,12'd4040};   
    1942 : result_out = {1'b1,12'd4041};   
    1943 : result_out = {1'b1,12'd4042};   
    1944 : result_out = {1'b1,12'd4043};   
    1945 : result_out = {1'b1,12'd4044};   
    1946 : result_out = {1'b1,12'd4045};   
    1947 : result_out = {1'b1,12'd4046};   
    1948 : result_out = {1'b1,12'd4047};   
    1949 : result_out = {1'b1,12'd4048};   
    1950 : result_out = {1'b1,12'd4049};   
    1951 : result_out = {1'b1,12'd4050};   
    1952 : result_out = {1'b1,12'd4051};   
    1953 : result_out = {1'b1,12'd4052};   
    1954 : result_out = {1'b1,12'd4052};   
    1955 : result_out = {1'b1,12'd4053};   
    1956 : result_out = {1'b1,12'd4054};   
    1957 : result_out = {1'b1,12'd4055};   
    1958 : result_out = {1'b1,12'd4056};   
    1959 : result_out = {1'b1,12'd4057};   
    1960 : result_out = {1'b1,12'd4058};   
    1961 : result_out = {1'b1,12'd4059};   
    1962 : result_out = {1'b1,12'd4059};   
    1963 : result_out = {1'b1,12'd4060};   
    1964 : result_out = {1'b1,12'd4061};   
    1965 : result_out = {1'b1,12'd4062};   
    1966 : result_out = {1'b1,12'd4063};   
    1967 : result_out = {1'b1,12'd4063};   
    1968 : result_out = {1'b1,12'd4064};   
    1969 : result_out = {1'b1,12'd4065};   
    1970 : result_out = {1'b1,12'd4066};   
    1971 : result_out = {1'b1,12'd4066};   
    1972 : result_out = {1'b1,12'd4067};   
    1973 : result_out = {1'b1,12'd4068};   
    1974 : result_out = {1'b1,12'd4069};   
    1975 : result_out = {1'b1,12'd4069};   
    1976 : result_out = {1'b1,12'd4070};   
    1977 : result_out = {1'b1,12'd4071};   
    1978 : result_out = {1'b1,12'd4071};   
    1979 : result_out = {1'b1,12'd4072};   
    1980 : result_out = {1'b1,12'd4073};   
    1981 : result_out = {1'b1,12'd4073};   
    1982 : result_out = {1'b1,12'd4074};   
    1983 : result_out = {1'b1,12'd4075};   
    1984 : result_out = {1'b1,12'd4075};   
    1985 : result_out = {1'b1,12'd4076};   
    1986 : result_out = {1'b1,12'd4076};   
    1987 : result_out = {1'b1,12'd4077};   
    1988 : result_out = {1'b1,12'd4078};   
    1989 : result_out = {1'b1,12'd4078};   
    1990 : result_out = {1'b1,12'd4079};   
    1991 : result_out = {1'b1,12'd4079};   
    1992 : result_out = {1'b1,12'd4080};   
    1993 : result_out = {1'b1,12'd4080};   
    1994 : result_out = {1'b1,12'd4081};   
    1995 : result_out = {1'b1,12'd4081};   
    1996 : result_out = {1'b1,12'd4082};   
    1997 : result_out = {1'b1,12'd4082};   
    1998 : result_out = {1'b1,12'd4083};   
    1999 : result_out = {1'b1,12'd4083};   
    2000 : result_out = {1'b1,12'd4084};   
    2001 : result_out = {1'b1,12'd4084};   
    2002 : result_out = {1'b1,12'd4085};   
    2003 : result_out = {1'b1,12'd4085};   
    2004 : result_out = {1'b1,12'd4086};   
    2005 : result_out = {1'b1,12'd4086};   
    2006 : result_out = {1'b1,12'd4087};   
    2007 : result_out = {1'b1,12'd4087};   
    2008 : result_out = {1'b1,12'd4087};   
    2009 : result_out = {1'b1,12'd4088};   
    2010 : result_out = {1'b1,12'd4088};   
    2011 : result_out = {1'b1,12'd4088};   
    2012 : result_out = {1'b1,12'd4089};   
    2013 : result_out = {1'b1,12'd4089};   
    2014 : result_out = {1'b1,12'd4089};   
    2015 : result_out = {1'b1,12'd4090};   
    2016 : result_out = {1'b1,12'd4090};   
    2017 : result_out = {1'b1,12'd4090};   
    2018 : result_out = {1'b1,12'd4091};   
    2019 : result_out = {1'b1,12'd4091};   
    2020 : result_out = {1'b1,12'd4091};   
    2021 : result_out = {1'b1,12'd4091};   
    2022 : result_out = {1'b1,12'd4092};   
    2023 : result_out = {1'b1,12'd4092};   
    2024 : result_out = {1'b1,12'd4092};   
    2025 : result_out = {1'b1,12'd4092};   
    2026 : result_out = {1'b1,12'd4093};   
    2027 : result_out = {1'b1,12'd4093};   
    2028 : result_out = {1'b1,12'd4093};   
    2029 : result_out = {1'b1,12'd4093};   
    2030 : result_out = {1'b1,12'd4093};   
    2031 : result_out = {1'b1,12'd4094};   
    2032 : result_out = {1'b1,12'd4094};   
    2033 : result_out = {1'b1,12'd4094};   
    2034 : result_out = {1'b1,12'd4094};   
    2035 : result_out = {1'b1,12'd4094};   
    2036 : result_out = {1'b1,12'd4094};   
    2037 : result_out = {1'b1,12'd4094};   
    2038 : result_out = {1'b1,12'd4095};   
    2039 : result_out = {1'b1,12'd4095};   
    2040 : result_out = {1'b1,12'd4095};   
    2041 : result_out = {1'b1,12'd4095};   
    2042 : result_out = {1'b1,12'd4095};   
    2043 : result_out = {1'b1,12'd4095};   
    2044 : result_out = {1'b1,12'd4095};   
    2045 : result_out = {1'b1,12'd4095};   
    2046 : result_out = {1'b1,12'd4095};   
    2047 : result_out = {1'b1,12'd4095};   
    2048 : result_out = {1'b1,12'd4095};   
    default: result_out = {1'b0,x_in}; // Default case
    endcase
end

endmodule



