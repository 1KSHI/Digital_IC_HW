module Divder12(
    input [23:0] x_in,
    input [23:0] y_in,
    output [23:0] result_out
);

assign result_out = x_in/y_in;

endmodule
